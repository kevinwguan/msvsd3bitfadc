magic
tech sky130A
timestamp 1676772270
<< nwell >>
rect 10 320 670 670
<< nmos >>
rect 120 90 140 260
rect 200 90 220 260
rect 280 90 300 260
rect 360 90 380 260
rect 440 90 460 260
rect 520 90 540 260
<< pmos >>
rect 120 380 140 550
rect 200 380 220 550
rect 280 380 300 550
rect 360 380 380 550
rect 440 380 460 550
rect 520 380 540 550
<< ndiff >>
rect 60 220 70 260
rect 110 220 120 260
rect 60 90 120 220
rect 140 200 200 260
rect 140 160 150 200
rect 190 160 200 200
rect 140 90 200 160
rect 220 220 230 260
rect 270 220 280 260
rect 220 90 280 220
rect 300 90 360 260
rect 380 130 440 260
rect 380 90 390 130
rect 430 90 440 130
rect 460 200 520 260
rect 460 160 470 200
rect 510 160 520 200
rect 460 90 520 160
rect 540 130 600 260
rect 540 90 550 130
rect 590 90 600 130
<< pdiff >>
rect 60 510 70 550
rect 110 510 120 550
rect 60 380 120 510
rect 140 380 200 550
rect 220 510 230 550
rect 270 510 280 550
rect 220 380 280 510
rect 300 420 360 550
rect 300 380 310 420
rect 350 380 360 420
rect 380 510 390 550
rect 430 510 440 550
rect 380 380 440 510
rect 460 380 520 550
rect 540 510 550 550
rect 590 510 600 550
rect 540 380 600 510
<< ndiffc >>
rect 70 220 110 260
rect 150 160 190 200
rect 230 220 270 260
rect 390 90 430 130
rect 470 160 510 200
rect 550 90 590 130
<< pdiffc >>
rect 70 510 110 550
rect 230 510 270 550
rect 310 380 350 420
rect 390 510 430 550
rect 550 510 590 550
<< psubdiffcont >>
rect 40 10 80 40
rect 120 10 160 40
rect 200 10 240 40
rect 280 10 320 40
rect 360 10 400 40
rect 440 10 480 40
rect 520 10 560 40
rect 600 10 640 40
<< nsubdiffcont >>
rect 40 600 80 640
rect 120 600 160 640
rect 200 600 240 640
rect 280 600 320 640
rect 360 600 400 640
rect 440 600 480 640
rect 520 600 560 640
rect 600 600 640 640
<< poly >>
rect 120 550 140 580
rect 200 550 220 580
rect 280 550 300 580
rect 360 550 380 580
rect 440 550 460 580
rect 520 550 540 580
rect 120 260 140 380
rect 200 260 220 380
rect 280 260 300 380
rect 360 260 380 380
rect 440 260 460 380
rect 520 260 540 380
rect 120 60 140 90
rect 200 60 220 90
rect 280 60 300 90
rect 360 60 380 90
rect 440 60 460 90
rect 520 60 540 90
<< metal1 >>
rect 10 600 40 640
rect 80 600 120 640
rect 160 600 200 640
rect 240 600 280 640
rect 320 600 360 640
rect 400 600 440 640
rect 480 600 520 640
rect 560 600 600 640
rect 640 600 660 640
rect 70 550 110 600
rect 550 550 580 600
rect 270 520 390 550
rect 310 320 340 380
rect 70 290 340 320
rect 70 260 100 290
rect 230 260 260 290
rect 190 160 470 190
rect 390 40 430 90
rect 550 40 590 90
rect 10 10 40 40
rect 80 10 120 40
rect 160 10 200 40
rect 240 10 280 40
rect 320 10 360 40
rect 400 10 440 40
rect 480 10 520 40
rect 560 10 600 40
rect 640 10 660 40
<< labels >>
rlabel pdiffc 550 510 590 550 1 vdd
port 1 n
rlabel pdiffc 70 510 110 550 1 vdd
rlabel ndiffc 550 90 590 130 1 gnd
port 3 n
rlabel ndiffc 390 90 430 130 1 gnd
rlabel pdiffc 310 380 350 420 1 out
rlabel ndiffc 230 220 270 260 1 out
rlabel ndiffc 70 220 110 260 1 out
port 2 n
rlabel poly 120 260 140 380 1 a
port 4 n
rlabel poly 520 260 540 380 1 b
port 9 n
rlabel poly 200 260 220 380 1 c
port 5 n
rlabel poly 440 260 460 380 1 d
port 8 n
rlabel poly 280 260 300 380 1 e
port 6 n
rlabel poly 360 260 380 380 1 f
port 7 n
<< end >>
