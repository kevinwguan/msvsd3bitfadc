* NGSPICE file created from fn_postlayout.ext - technology: sky130A

.subckt fn_postlayout vdd out gnd a c e f d b
X0 a_280_760# a vdd w_20_640# sky130_fd_pr__pfet_01v8 ad=1.02e+12p pd=4.6e+06u as=2.04e+12p ps=9.2e+06u w=1.7e+06u l=200000u
X1 a_760_760# f out w_20_640# sky130_fd_pr__pfet_01v8 ad=1.02e+12p pd=4.6e+06u as=1.02e+12p ps=4.6e+06u w=1.7e+06u l=200000u
X2 a_600_180# e out a_80_20# sky130_fd_pr__nfet_01v8 ad=1.02e+12p pd=4.6e+06u as=2.04e+12p ps=9.2e+06u w=1.7e+06u l=200000u
X3 gnd b a_920_180# a_80_20# sky130_fd_pr__nfet_01v8 ad=2.04e+12p pd=9.2e+06u as=1.02e+12p ps=4.6e+06u w=1.7e+06u l=200000u
X4 a_920_760# d a_760_760# w_20_640# sky130_fd_pr__pfet_01v8 ad=1.02e+12p pd=4.6e+06u as=0p ps=0u w=1.7e+06u l=200000u
X5 a_440_760# c a_280_760# w_20_640# sky130_fd_pr__pfet_01v8 ad=1.02e+12p pd=4.6e+06u as=0p ps=0u w=1.7e+06u l=200000u
X6 a_280_180# a out a_80_20# sky130_fd_pr__nfet_01v8 ad=1.02e+12p pd=4.6e+06u as=0p ps=0u w=1.7e+06u l=200000u
X7 gnd f a_600_180# a_80_20# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.7e+06u l=200000u
X8 out e a_440_760# w_20_640# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.7e+06u l=200000u
X9 a_920_180# d gnd a_80_20# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.7e+06u l=200000u
X10 vdd b a_920_760# w_20_640# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.7e+06u l=200000u
X11 out c a_280_180# a_80_20# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.7e+06u l=200000u
.ends

