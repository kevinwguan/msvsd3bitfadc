* NGSPICE file created from SECTION7.ext - technology: sky130A

.subckt SECTION7 vdd gnd out 1 2 3 4 5 6
X0 out 2 a_663_2352# vdd sky130_fd_pr__pfet_01v8 ad=2.94e+11p pd=2.66e+06u as=8.505e+11p ps=7.92e+06u w=1.05e+06u l=150000u
X1 a_230_2352# 3 a_1262_2352# vdd sky130_fd_pr__pfet_01v8 ad=8.505e+11p pd=7.92e+06u as=8.505e+11p ps=7.92e+06u w=1.05e+06u l=150000u
X2 a_230_2352# 1 a_147_2352# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.565e+11p ps=5.26e+06u w=1.05e+06u l=150000u
X3 a_663_2352# 2 out vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X4 a_1695_462# 4 a_663_462# gnd sky130_fd_pr__nfet_01v8 ad=8.505e+11p pd=7.92e+06u as=8.505e+11p ps=7.92e+06u w=1.05e+06u l=150000u
X5 a_1262_462# 5 a_2294_462# gnd sky130_fd_pr__nfet_01v8 ad=8.505e+11p pd=7.92e+06u as=8.505e+11p ps=7.92e+06u w=1.05e+06u l=150000u
X6 a_147_2352# 1 a_230_2352# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X7 a_663_2352# 4 a_1695_2352# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.505e+11p ps=7.92e+06u w=1.05e+06u l=150000u
X8 out 2 a_663_462# gnd sky130_fd_pr__nfet_01v8 ad=2.94e+11p pd=2.66e+06u as=0p ps=0u w=1.05e+06u l=150000u
X9 a_1695_462# 6 a_2294_462# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X10 a_1262_2352# 3 a_230_2352# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X11 a_1695_2352# 4 a_663_2352# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X12 a_663_462# 2 out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X13 a_2294_462# 6 a_1695_462# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X14 a_1262_462# 3 a_230_462# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.505e+11p ps=7.92e+06u w=1.05e+06u l=150000u
X15 a_2294_2352# 5 a_1262_2352# vdd sky130_fd_pr__pfet_01v8 ad=8.505e+11p pd=7.92e+06u as=0p ps=0u w=1.05e+06u l=150000u
X16 a_2294_2352# 6 a_1695_2352# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X17 a_1262_2352# 5 a_2294_2352# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X18 a_230_462# 3 a_1262_462# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X19 a_230_462# 1 a_147_462# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.565e+11p ps=5.26e+06u w=1.05e+06u l=150000u
X20 a_147_462# 1 a_230_462# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X21 a_663_462# 4 a_1695_462# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X22 a_1695_2352# 6 a_2294_2352# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X23 a_2294_462# 5 a_1262_462# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
.ends

