MACRO ADC_FINAL
  ORIGIN 0 0 ;
  FOREIGN ADC_FINAL 0 0 ;
  SIZE 16.34 BY 15.12 ;
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.15 7.82 1.43 8.98 ;
      LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
      LAYER M2 ;
        RECT 5.42 7 10.06 7.28 ;
      LAYER M3 ;
        RECT 1.15 7.56 1.43 7.98 ;
      LAYER M2 ;
        RECT 1.29 7.42 3.01 7.7 ;
      LAYER M1 ;
        RECT 2.885 7.56 3.135 7.98 ;
      LAYER M2 ;
        RECT 2.85 7.84 3.17 8.12 ;
      LAYER M2 ;
        RECT 3.87 7.84 4.73 8.12 ;
      LAYER M1 ;
        RECT 4.605 7.14 4.855 7.98 ;
      LAYER M2 ;
        RECT 4.73 7 5.59 7.28 ;
    END
  END VOUT
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 8.03 0.68 8.31 6.88 ;
      LAYER M3 ;
        RECT 14.05 0.68 14.33 6.46 ;
      LAYER M3 ;
        RECT 8.03 1.075 8.31 1.445 ;
      LAYER M2 ;
        RECT 8.17 1.12 14.19 1.4 ;
      LAYER M3 ;
        RECT 14.05 1.075 14.33 1.445 ;
      LAYER M2 ;
        RECT 8.86 14.14 10.92 14.42 ;
      LAYER M2 ;
        RECT 13.16 14.14 15.22 14.42 ;
      LAYER M3 ;
        RECT 8.03 6.72 8.31 14.28 ;
      LAYER M2 ;
        RECT 8.17 14.14 9.03 14.42 ;
      LAYER M2 ;
        RECT 10.75 14.14 13.33 14.42 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 2.01 0.68 2.29 6.46 ;
      LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
      LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
      LAYER M2 ;
        RECT 1.12 14.14 2.32 14.42 ;
      LAYER M3 ;
        RECT 2.01 6.115 2.29 6.485 ;
      LAYER M4 ;
        RECT 2.15 5.9 4.3 6.7 ;
      LAYER M3 ;
        RECT 4.16 6.3 4.44 8.4 ;
      LAYER M3 ;
        RECT 4.16 8.635 4.44 9.005 ;
      LAYER M2 ;
        RECT 4.3 8.68 6.02 8.96 ;
      LAYER M3 ;
        RECT 5.88 8.635 6.16 9.005 ;
      LAYER M3 ;
        RECT 4.16 13.675 4.44 14.045 ;
      LAYER M2 ;
        RECT 2.15 13.72 4.3 14 ;
      LAYER M1 ;
        RECT 2.025 13.86 2.275 14.28 ;
      LAYER M2 ;
        RECT 1.99 14.14 2.31 14.42 ;
    END
  END VSS
  PIN VPOS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 13.16 12.04 15.22 12.32 ;
    END
  END VPOS
  OBS 
  LAYER M2 ;
        RECT 5.42 2.8 10.06 3.08 ;
  LAYER M3 ;
        RECT 13.19 2.78 13.47 7.3 ;
  LAYER M2 ;
        RECT 9.89 2.8 11.61 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.94 11.75 3.36 ;
  LAYER M2 ;
        RECT 11.61 3.22 13.33 3.5 ;
  LAYER M3 ;
        RECT 13.19 3.175 13.47 3.545 ;
  LAYER M3 ;
        RECT 6.31 7.82 6.59 12.34 ;
  LAYER M2 ;
        RECT 8.86 12.04 10.92 12.32 ;
  LAYER M2 ;
        RECT 6.29 2.8 6.61 3.08 ;
  LAYER M3 ;
        RECT 6.31 2.94 6.59 7.98 ;
  LAYER M3 ;
        RECT 6.31 11.575 6.59 11.945 ;
  LAYER M2 ;
        RECT 6.45 11.62 8.6 11.9 ;
  LAYER M1 ;
        RECT 8.475 11.76 8.725 12.18 ;
  LAYER M2 ;
        RECT 8.6 12.04 9.03 12.32 ;
  LAYER M2 ;
        RECT 6.29 2.8 6.61 3.08 ;
  LAYER M3 ;
        RECT 6.31 2.78 6.59 3.1 ;
  LAYER M2 ;
        RECT 6.29 2.8 6.61 3.08 ;
  LAYER M3 ;
        RECT 6.31 2.78 6.59 3.1 ;
  LAYER M1 ;
        RECT 8.475 11.675 8.725 11.845 ;
  LAYER M2 ;
        RECT 8.43 11.62 8.77 11.9 ;
  LAYER M1 ;
        RECT 8.475 12.095 8.725 12.265 ;
  LAYER M2 ;
        RECT 8.43 12.04 8.77 12.32 ;
  LAYER M2 ;
        RECT 6.29 2.8 6.61 3.08 ;
  LAYER M3 ;
        RECT 6.31 2.78 6.59 3.1 ;
  LAYER M2 ;
        RECT 6.29 11.62 6.61 11.9 ;
  LAYER M3 ;
        RECT 6.31 11.6 6.59 11.92 ;
  LAYER M1 ;
        RECT 8.475 11.675 8.725 11.845 ;
  LAYER M2 ;
        RECT 8.43 11.62 8.77 11.9 ;
  LAYER M1 ;
        RECT 8.475 12.095 8.725 12.265 ;
  LAYER M2 ;
        RECT 8.43 12.04 8.77 12.32 ;
  LAYER M2 ;
        RECT 6.29 2.8 6.61 3.08 ;
  LAYER M3 ;
        RECT 6.31 2.78 6.59 3.1 ;
  LAYER M2 ;
        RECT 6.29 11.62 6.61 11.9 ;
  LAYER M3 ;
        RECT 6.31 11.6 6.59 11.92 ;
  LAYER M2 ;
        RECT 8.43 8.26 11.35 8.54 ;
  LAYER M2 ;
        RECT 12.73 8.26 15.65 8.54 ;
  LAYER M2 ;
        RECT 12.3 6.58 15.22 6.86 ;
  LAYER M2 ;
        RECT 11.18 8.26 12.9 8.54 ;
  LAYER M2 ;
        RECT 12.31 8.26 12.63 8.54 ;
  LAYER M3 ;
        RECT 12.33 6.72 12.61 8.4 ;
  LAYER M2 ;
        RECT 12.31 6.58 12.63 6.86 ;
  LAYER M2 ;
        RECT 12.31 6.58 12.63 6.86 ;
  LAYER M3 ;
        RECT 12.33 6.56 12.61 6.88 ;
  LAYER M2 ;
        RECT 12.31 8.26 12.63 8.54 ;
  LAYER M3 ;
        RECT 12.33 8.24 12.61 8.56 ;
  LAYER M2 ;
        RECT 12.31 6.58 12.63 6.86 ;
  LAYER M3 ;
        RECT 12.33 6.56 12.61 6.88 ;
  LAYER M2 ;
        RECT 12.31 8.26 12.63 8.54 ;
  LAYER M3 ;
        RECT 12.33 8.24 12.61 8.56 ;
  LAYER M3 ;
        RECT 2.87 2.78 3.15 7.3 ;
  LAYER M2 ;
        RECT 8.86 7.84 10.92 8.12 ;
  LAYER M3 ;
        RECT 2.87 7.14 3.15 7.56 ;
  LAYER M4 ;
        RECT 3.01 7.16 8.6 7.96 ;
  LAYER M3 ;
        RECT 8.46 7.56 8.74 7.98 ;
  LAYER M2 ;
        RECT 8.6 7.84 9.03 8.12 ;
  LAYER M2 ;
        RECT 8.44 7.84 8.76 8.12 ;
  LAYER M3 ;
        RECT 8.46 7.82 8.74 8.14 ;
  LAYER M3 ;
        RECT 2.87 7.375 3.15 7.745 ;
  LAYER M4 ;
        RECT 2.845 7.16 3.175 7.96 ;
  LAYER M3 ;
        RECT 8.46 7.375 8.74 7.745 ;
  LAYER M4 ;
        RECT 8.435 7.16 8.765 7.96 ;
  LAYER M2 ;
        RECT 8.44 7.84 8.76 8.12 ;
  LAYER M3 ;
        RECT 8.46 7.82 8.74 8.14 ;
  LAYER M3 ;
        RECT 2.87 7.375 3.15 7.745 ;
  LAYER M4 ;
        RECT 2.845 7.16 3.175 7.96 ;
  LAYER M3 ;
        RECT 8.46 7.375 8.74 7.745 ;
  LAYER M4 ;
        RECT 8.435 7.16 8.765 7.96 ;
  LAYER M2 ;
        RECT 1.98 6.58 3.18 6.86 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M2 ;
        RECT 13.16 7.84 15.22 8.12 ;
  LAYER M2 ;
        RECT 1.72 6.58 2.15 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.72 1.86 12.18 ;
  LAYER M2 ;
        RECT 1.56 12.04 1.88 12.32 ;
  LAYER M2 ;
        RECT 2.15 12.04 3.01 12.32 ;
  LAYER M2 ;
        RECT 3.01 6.58 4.3 6.86 ;
  LAYER M1 ;
        RECT 4.175 6.72 4.425 7.56 ;
  LAYER M2 ;
        RECT 4.3 7.42 12.47 7.7 ;
  LAYER M1 ;
        RECT 12.345 7.56 12.595 7.98 ;
  LAYER M2 ;
        RECT 12.47 7.84 13.33 8.12 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 12.04 1.88 12.32 ;
  LAYER M3 ;
        RECT 1.58 12.02 1.86 12.34 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 12.04 1.88 12.32 ;
  LAYER M3 ;
        RECT 1.58 12.02 1.86 12.34 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 12.04 1.88 12.32 ;
  LAYER M3 ;
        RECT 1.58 12.02 1.86 12.34 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 12.04 1.88 12.32 ;
  LAYER M3 ;
        RECT 1.58 12.02 1.86 12.34 ;
  LAYER M1 ;
        RECT 4.175 6.635 4.425 6.805 ;
  LAYER M2 ;
        RECT 4.13 6.58 4.47 6.86 ;
  LAYER M1 ;
        RECT 4.175 7.475 4.425 7.645 ;
  LAYER M2 ;
        RECT 4.13 7.42 4.47 7.7 ;
  LAYER M1 ;
        RECT 12.345 7.475 12.595 7.645 ;
  LAYER M2 ;
        RECT 12.3 7.42 12.64 7.7 ;
  LAYER M1 ;
        RECT 12.345 7.895 12.595 8.065 ;
  LAYER M2 ;
        RECT 12.3 7.84 12.64 8.12 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 12.04 1.88 12.32 ;
  LAYER M3 ;
        RECT 1.58 12.02 1.86 12.34 ;
  LAYER M1 ;
        RECT 4.175 6.635 4.425 6.805 ;
  LAYER M2 ;
        RECT 4.13 6.58 4.47 6.86 ;
  LAYER M1 ;
        RECT 4.175 7.475 4.425 7.645 ;
  LAYER M2 ;
        RECT 4.13 7.42 4.47 7.7 ;
  LAYER M1 ;
        RECT 12.345 7.475 12.595 7.645 ;
  LAYER M2 ;
        RECT 12.3 7.42 12.64 7.7 ;
  LAYER M1 ;
        RECT 12.345 7.895 12.595 8.065 ;
  LAYER M2 ;
        RECT 12.3 7.84 12.64 8.12 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 12.04 1.88 12.32 ;
  LAYER M3 ;
        RECT 1.58 12.02 1.86 12.34 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M2 ;
        RECT 13.16 7 14.36 7.28 ;
  LAYER M2 ;
        RECT 12.3 2.8 15.22 3.08 ;
  LAYER M2 ;
        RECT 12.3 0.7 15.22 0.98 ;
  LAYER M2 ;
        RECT 11.87 6.16 15.65 6.44 ;
  LAYER M3 ;
        RECT 13.19 2.78 13.47 7.3 ;
  LAYER M2 ;
        RECT 12.3 6.58 15.22 6.86 ;
  LAYER M3 ;
        RECT 14.05 0.68 14.33 6.46 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M2 ;
        RECT 5.42 0.7 10.06 0.98 ;
  LAYER M2 ;
        RECT 4.99 6.58 10.49 6.86 ;
  LAYER M2 ;
        RECT 5.42 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 5.42 2.8 10.06 3.08 ;
  LAYER M3 ;
        RECT 8.03 0.68 8.31 6.88 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 2.84 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 1.98 2.8 3.18 3.08 ;
  LAYER M2 ;
        RECT 1.98 0.7 3.18 0.98 ;
  LAYER M2 ;
        RECT 1.55 6.16 3.61 6.44 ;
  LAYER M3 ;
        RECT 2.87 2.78 3.15 7.3 ;
  LAYER M2 ;
        RECT 1.98 6.58 3.18 6.86 ;
  LAYER M3 ;
        RECT 2.01 0.68 2.29 6.46 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M3 ;
        RECT 6.31 7.82 6.59 12.34 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 1.12 14.14 2.32 14.42 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M3 ;
        RECT 1.15 7.82 1.43 8.98 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 11.425 ;
  LAYER M1 ;
        RECT 10.625 11.675 10.875 12.685 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 14.785 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M2 ;
        RECT 8.86 14.14 10.92 14.42 ;
  LAYER M2 ;
        RECT 8.86 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 8.86 12.04 10.92 12.32 ;
  LAYER M2 ;
        RECT 8.43 8.26 11.35 8.54 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 11.425 ;
  LAYER M1 ;
        RECT 14.925 11.675 15.175 12.685 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 14.785 ;
  LAYER M1 ;
        RECT 15.355 7.895 15.605 11.425 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 14.785 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 11.425 ;
  LAYER M1 ;
        RECT 13.205 11.675 13.455 12.685 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 14.785 ;
  LAYER M1 ;
        RECT 12.775 7.895 13.025 11.425 ;
  LAYER M2 ;
        RECT 13.16 14.14 15.22 14.42 ;
  LAYER M2 ;
        RECT 13.16 7.84 15.22 8.12 ;
  LAYER M2 ;
        RECT 13.16 12.04 15.22 12.32 ;
  LAYER M2 ;
        RECT 12.73 8.26 15.65 8.54 ;
  END 
END ADC_FINAL
