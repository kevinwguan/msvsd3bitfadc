.subckt section7 vdd out gnd a c e f d b
M0 10 c 9 a_8_0# sky130_fd_pr__nfet_01v8 w=10.5e-7 l=150e-9
M1 4 e 3 15 sky130_fd_pr__pfet_01v8 w=10.5e-7 l=150e-9
M2 3 c 2 15 sky130_fd_pr__pfet_01v8 w=10.5e-7 l=150e-9
M3 13 d 12 a_8_0# sky130_fd_pr__nfet_01v8 w=10.5e-7 l=150e-9
M4 12 f 11 a_8_0# sky130_fd_pr__nfet_01v8 w=10.5e-7 l=150e-9
M5 9 a 8 a_8_0# sky130_fd_pr__nfet_01v8 w=10.5e-7 l=150e-9
M6 14 b 13 a_8_0# sky130_fd_pr__nfet_01v8 w=10.5e-7 l=150e-9
M7 6 d 5 15 sky130_fd_pr__pfet_01v8 w=10.5e-7 l=150e-9
M8 5 f 4 15 sky130_fd_pr__pfet_01v8 w=10.5e-7 l=150e-9
M9 2 a 1 15 sky130_fd_pr__pfet_01v8 w=10.5e-7 l=150e-9
M10 7 b 6 15 sky130_fd_pr__pfet_01v8 w=10.5e-7 l=150e-9
M11 11 e 10 a_8_0# sky130_fd_pr__nfet_01v8 w=10.5e-7 l=150e-9
.ends section7

