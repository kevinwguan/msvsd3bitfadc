MACRO STAGE2_INV_91993238
  ORIGIN 0 0 ;
  FOREIGN STAGE2_INV_91993238 0 0 ;
  SIZE 5.16 BY 15.12 ;
  PIN VI
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
      LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
      LAYER M2 ;
        RECT 4.57 12.04 4.89 12.32 ;
      LAYER M3 ;
        RECT 4.59 2.94 4.87 12.18 ;
      LAYER M2 ;
        RECT 4.57 2.8 4.89 3.08 ;
    END
  END VI
  PIN SN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
      LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
      LAYER M3 ;
        RECT 3.3 6.115 3.58 6.485 ;
      LAYER M2 ;
        RECT 1.72 6.16 3.44 6.44 ;
      LAYER M3 ;
        RECT 1.58 6.115 1.86 6.485 ;
    END
  END SN
  PIN VO
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
      LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
      LAYER M2 ;
        RECT 0.27 7.84 0.59 8.12 ;
      LAYER M1 ;
        RECT 0.305 7.14 0.555 7.98 ;
      LAYER M2 ;
        RECT 0.27 7 0.59 7.28 ;
    END
  END VO
  PIN SP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
      LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
      LAYER M3 ;
        RECT 3.3 13.675 3.58 14.045 ;
      LAYER M2 ;
        RECT 1.72 13.72 3.44 14 ;
      LAYER M3 ;
        RECT 1.58 13.675 1.86 14.045 ;
    END
  END SP
  OBS 
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M2 ;
        RECT 1.29 12.04 3.01 12.32 ;
  LAYER M1 ;
        RECT 2.885 7.98 3.135 12.18 ;
  LAYER M2 ;
        RECT 3.01 7.84 3.87 8.12 ;
  LAYER M2 ;
        RECT 4.57 7.84 4.89 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.14 4.855 7.98 ;
  LAYER M2 ;
        RECT 4.57 7 4.89 7.28 ;
  LAYER M1 ;
        RECT 2.885 2.94 3.135 7.98 ;
  LAYER M2 ;
        RECT 1.29 2.8 3.01 3.08 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 2.885 2.855 3.135 3.025 ;
  LAYER M2 ;
        RECT 2.84 2.8 3.18 3.08 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 2.885 2.855 3.135 3.025 ;
  LAYER M2 ;
        RECT 2.84 2.8 3.18 3.08 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  END 
END STAGE2_INV_91993238
