MACRO PMOS_S_2470631_X8_Y3
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN PMOS_S_2470631_X8_Y3 0 0 ;
  SIZE 8600 BY 19320 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 3730 260 4010 12340 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 4160 4460 4440 16540 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 4590 680 4870 18640 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 18985 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 18985 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M1 ;
      RECT 2885 335 3135 3865 ;
    LAYER M1 ;
      RECT 2885 4115 3135 5125 ;
    LAYER M1 ;
      RECT 2885 6215 3135 9745 ;
    LAYER M1 ;
      RECT 2885 9995 3135 11005 ;
    LAYER M1 ;
      RECT 2885 12095 3135 15625 ;
    LAYER M1 ;
      RECT 2885 15875 3135 16885 ;
    LAYER M1 ;
      RECT 2885 17975 3135 18985 ;
    LAYER M1 ;
      RECT 3315 335 3565 3865 ;
    LAYER M1 ;
      RECT 3315 6215 3565 9745 ;
    LAYER M1 ;
      RECT 3315 12095 3565 15625 ;
    LAYER M1 ;
      RECT 3745 335 3995 3865 ;
    LAYER M1 ;
      RECT 3745 4115 3995 5125 ;
    LAYER M1 ;
      RECT 3745 6215 3995 9745 ;
    LAYER M1 ;
      RECT 3745 9995 3995 11005 ;
    LAYER M1 ;
      RECT 3745 12095 3995 15625 ;
    LAYER M1 ;
      RECT 3745 15875 3995 16885 ;
    LAYER M1 ;
      RECT 3745 17975 3995 18985 ;
    LAYER M1 ;
      RECT 4175 335 4425 3865 ;
    LAYER M1 ;
      RECT 4175 6215 4425 9745 ;
    LAYER M1 ;
      RECT 4175 12095 4425 15625 ;
    LAYER M1 ;
      RECT 4605 335 4855 3865 ;
    LAYER M1 ;
      RECT 4605 4115 4855 5125 ;
    LAYER M1 ;
      RECT 4605 6215 4855 9745 ;
    LAYER M1 ;
      RECT 4605 9995 4855 11005 ;
    LAYER M1 ;
      RECT 4605 12095 4855 15625 ;
    LAYER M1 ;
      RECT 4605 15875 4855 16885 ;
    LAYER M1 ;
      RECT 4605 17975 4855 18985 ;
    LAYER M1 ;
      RECT 5035 335 5285 3865 ;
    LAYER M1 ;
      RECT 5035 6215 5285 9745 ;
    LAYER M1 ;
      RECT 5035 12095 5285 15625 ;
    LAYER M1 ;
      RECT 5465 335 5715 3865 ;
    LAYER M1 ;
      RECT 5465 4115 5715 5125 ;
    LAYER M1 ;
      RECT 5465 6215 5715 9745 ;
    LAYER M1 ;
      RECT 5465 9995 5715 11005 ;
    LAYER M1 ;
      RECT 5465 12095 5715 15625 ;
    LAYER M1 ;
      RECT 5465 15875 5715 16885 ;
    LAYER M1 ;
      RECT 5465 17975 5715 18985 ;
    LAYER M1 ;
      RECT 5895 335 6145 3865 ;
    LAYER M1 ;
      RECT 5895 6215 6145 9745 ;
    LAYER M1 ;
      RECT 5895 12095 6145 15625 ;
    LAYER M1 ;
      RECT 6325 335 6575 3865 ;
    LAYER M1 ;
      RECT 6325 4115 6575 5125 ;
    LAYER M1 ;
      RECT 6325 6215 6575 9745 ;
    LAYER M1 ;
      RECT 6325 9995 6575 11005 ;
    LAYER M1 ;
      RECT 6325 12095 6575 15625 ;
    LAYER M1 ;
      RECT 6325 15875 6575 16885 ;
    LAYER M1 ;
      RECT 6325 17975 6575 18985 ;
    LAYER M1 ;
      RECT 6755 335 7005 3865 ;
    LAYER M1 ;
      RECT 6755 6215 7005 9745 ;
    LAYER M1 ;
      RECT 6755 12095 7005 15625 ;
    LAYER M1 ;
      RECT 7185 335 7435 3865 ;
    LAYER M1 ;
      RECT 7185 4115 7435 5125 ;
    LAYER M1 ;
      RECT 7185 6215 7435 9745 ;
    LAYER M1 ;
      RECT 7185 9995 7435 11005 ;
    LAYER M1 ;
      RECT 7185 12095 7435 15625 ;
    LAYER M1 ;
      RECT 7185 15875 7435 16885 ;
    LAYER M1 ;
      RECT 7185 17975 7435 18985 ;
    LAYER M1 ;
      RECT 7615 335 7865 3865 ;
    LAYER M1 ;
      RECT 7615 6215 7865 9745 ;
    LAYER M1 ;
      RECT 7615 12095 7865 15625 ;
    LAYER M2 ;
      RECT 1120 280 7480 560 ;
    LAYER M2 ;
      RECT 1120 4480 7480 4760 ;
    LAYER M2 ;
      RECT 690 700 7910 980 ;
    LAYER M2 ;
      RECT 1120 6160 7480 6440 ;
    LAYER M2 ;
      RECT 1120 10360 7480 10640 ;
    LAYER M2 ;
      RECT 690 6580 7910 6860 ;
    LAYER M2 ;
      RECT 1120 12040 7480 12320 ;
    LAYER M2 ;
      RECT 1120 16240 7480 16520 ;
    LAYER M2 ;
      RECT 690 12460 7910 12740 ;
    LAYER M2 ;
      RECT 1120 18340 7480 18620 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 18395 1375 18565 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 18395 2235 18565 ;
    LAYER V1 ;
      RECT 2925 335 3095 505 ;
    LAYER V1 ;
      RECT 2925 4535 3095 4705 ;
    LAYER V1 ;
      RECT 2925 6215 3095 6385 ;
    LAYER V1 ;
      RECT 2925 10415 3095 10585 ;
    LAYER V1 ;
      RECT 2925 12095 3095 12265 ;
    LAYER V1 ;
      RECT 2925 16295 3095 16465 ;
    LAYER V1 ;
      RECT 2925 18395 3095 18565 ;
    LAYER V1 ;
      RECT 3785 335 3955 505 ;
    LAYER V1 ;
      RECT 3785 4535 3955 4705 ;
    LAYER V1 ;
      RECT 3785 6215 3955 6385 ;
    LAYER V1 ;
      RECT 3785 10415 3955 10585 ;
    LAYER V1 ;
      RECT 3785 12095 3955 12265 ;
    LAYER V1 ;
      RECT 3785 16295 3955 16465 ;
    LAYER V1 ;
      RECT 3785 18395 3955 18565 ;
    LAYER V1 ;
      RECT 4645 335 4815 505 ;
    LAYER V1 ;
      RECT 4645 4535 4815 4705 ;
    LAYER V1 ;
      RECT 4645 6215 4815 6385 ;
    LAYER V1 ;
      RECT 4645 10415 4815 10585 ;
    LAYER V1 ;
      RECT 4645 12095 4815 12265 ;
    LAYER V1 ;
      RECT 4645 16295 4815 16465 ;
    LAYER V1 ;
      RECT 4645 18395 4815 18565 ;
    LAYER V1 ;
      RECT 5505 335 5675 505 ;
    LAYER V1 ;
      RECT 5505 4535 5675 4705 ;
    LAYER V1 ;
      RECT 5505 6215 5675 6385 ;
    LAYER V1 ;
      RECT 5505 10415 5675 10585 ;
    LAYER V1 ;
      RECT 5505 12095 5675 12265 ;
    LAYER V1 ;
      RECT 5505 16295 5675 16465 ;
    LAYER V1 ;
      RECT 5505 18395 5675 18565 ;
    LAYER V1 ;
      RECT 6365 335 6535 505 ;
    LAYER V1 ;
      RECT 6365 4535 6535 4705 ;
    LAYER V1 ;
      RECT 6365 6215 6535 6385 ;
    LAYER V1 ;
      RECT 6365 10415 6535 10585 ;
    LAYER V1 ;
      RECT 6365 12095 6535 12265 ;
    LAYER V1 ;
      RECT 6365 16295 6535 16465 ;
    LAYER V1 ;
      RECT 6365 18395 6535 18565 ;
    LAYER V1 ;
      RECT 7225 335 7395 505 ;
    LAYER V1 ;
      RECT 7225 4535 7395 4705 ;
    LAYER V1 ;
      RECT 7225 6215 7395 6385 ;
    LAYER V1 ;
      RECT 7225 10415 7395 10585 ;
    LAYER V1 ;
      RECT 7225 12095 7395 12265 ;
    LAYER V1 ;
      RECT 7225 16295 7395 16465 ;
    LAYER V1 ;
      RECT 7225 18395 7395 18565 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V1 ;
      RECT 3355 755 3525 925 ;
    LAYER V1 ;
      RECT 3355 6635 3525 6805 ;
    LAYER V1 ;
      RECT 3355 12515 3525 12685 ;
    LAYER V1 ;
      RECT 4215 755 4385 925 ;
    LAYER V1 ;
      RECT 4215 6635 4385 6805 ;
    LAYER V1 ;
      RECT 4215 12515 4385 12685 ;
    LAYER V1 ;
      RECT 5075 755 5245 925 ;
    LAYER V1 ;
      RECT 5075 6635 5245 6805 ;
    LAYER V1 ;
      RECT 5075 12515 5245 12685 ;
    LAYER V1 ;
      RECT 5935 755 6105 925 ;
    LAYER V1 ;
      RECT 5935 6635 6105 6805 ;
    LAYER V1 ;
      RECT 5935 12515 6105 12685 ;
    LAYER V1 ;
      RECT 6795 755 6965 925 ;
    LAYER V1 ;
      RECT 6795 6635 6965 6805 ;
    LAYER V1 ;
      RECT 6795 12515 6965 12685 ;
    LAYER V1 ;
      RECT 7655 755 7825 925 ;
    LAYER V1 ;
      RECT 7655 6635 7825 6805 ;
    LAYER V1 ;
      RECT 7655 12515 7825 12685 ;
    LAYER V2 ;
      RECT 3795 345 3945 495 ;
    LAYER V2 ;
      RECT 3795 6225 3945 6375 ;
    LAYER V2 ;
      RECT 3795 12105 3945 12255 ;
    LAYER V2 ;
      RECT 4225 4545 4375 4695 ;
    LAYER V2 ;
      RECT 4225 10425 4375 10575 ;
    LAYER V2 ;
      RECT 4225 16305 4375 16455 ;
    LAYER V2 ;
      RECT 4655 765 4805 915 ;
    LAYER V2 ;
      RECT 4655 6645 4805 6795 ;
    LAYER V2 ;
      RECT 4655 12525 4805 12675 ;
    LAYER V2 ;
      RECT 4655 18405 4805 18555 ;
  END
END PMOS_S_2470631_X8_Y3
