** sch_path: /home/kevin/Documents/Day1/inverter/xschem/inverter_tb.sch
**.subckt inverter_tb out in
*.opin out
*.opin in
x1 gate vdd vss vout inverter
V1 gate vss pwl(0 0 1000n 1.8)
.save i(v1)
V2 vdd vss 1.8
.save i(v2)
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.control
	tran 1n 1u
	plot v(gate) v(vout)
.endc
.save all


**** end user architecture code
**.ends

.include inverter.spice

.GLOBAL vss
.end
