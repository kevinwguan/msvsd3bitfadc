MACRO SECTION7
  ORIGIN 0 0 ;
  FOREIGN SECTION7 0 0 ;
  SIZE 15.48 BY 15.12 ;
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 6.28 4.48 7.48 4.76 ;
      LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
      LAYER M2 ;
        RECT 6.72 4.48 7.04 4.76 ;
      LAYER M1 ;
        RECT 6.755 4.62 7.005 10.5 ;
      LAYER M2 ;
        RECT 6.72 10.36 7.04 10.64 ;
    END
  END C
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 11.44 4.48 12.64 4.76 ;
      LAYER M2 ;
        RECT 11.44 10.36 12.64 10.64 ;
      LAYER M2 ;
        RECT 11.88 4.48 12.2 4.76 ;
      LAYER M1 ;
        RECT 11.915 4.62 12.165 10.5 ;
      LAYER M2 ;
        RECT 11.88 10.36 12.2 10.64 ;
    END
  END E
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8 4.48 9.2 4.76 ;
      LAYER M2 ;
        RECT 8 10.36 9.2 10.64 ;
      LAYER M2 ;
        RECT 8.01 4.48 8.33 4.76 ;
      LAYER M1 ;
        RECT 8.045 4.62 8.295 10.5 ;
      LAYER M2 ;
        RECT 8.01 10.36 8.33 10.64 ;
    END
  END D
  PIN F
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 13.16 4.48 14.36 4.76 ;
      LAYER M2 ;
        RECT 13.16 10.36 14.36 10.64 ;
      LAYER M2 ;
        RECT 13.17 4.48 13.49 4.76 ;
      LAYER M1 ;
        RECT 13.205 4.62 13.455 10.5 ;
      LAYER M2 ;
        RECT 13.17 10.36 13.49 10.64 ;
    END
  END F
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 4.48 2.32 4.76 ;
      LAYER M2 ;
        RECT 1.12 10.36 2.32 10.64 ;
      LAYER M2 ;
        RECT 1.56 4.48 1.88 4.76 ;
      LAYER M1 ;
        RECT 1.595 4.62 1.845 10.5 ;
      LAYER M2 ;
        RECT 1.56 10.36 1.88 10.64 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 2.84 4.48 4.04 4.76 ;
      LAYER M2 ;
        RECT 2.84 10.36 4.04 10.64 ;
      LAYER M2 ;
        RECT 2.85 4.48 3.17 4.76 ;
      LAYER M1 ;
        RECT 2.885 4.62 3.135 10.5 ;
      LAYER M2 ;
        RECT 2.85 10.36 3.17 10.64 ;
    END
  END B
  OBS 
  LAYER M2 ;
        RECT 1.12 6.58 2.32 6.86 ;
  LAYER M2 ;
        RECT 2.84 6.58 4.04 6.86 ;
  LAYER M2 ;
        RECT 6.28 6.58 7.48 6.86 ;
  LAYER M2 ;
        RECT 8 6.58 9.2 6.86 ;
  LAYER M2 ;
        RECT 11.44 6.58 12.64 6.86 ;
  LAYER M2 ;
        RECT 13.16 6.58 14.36 6.86 ;
  LAYER M2 ;
        RECT 2.15 6.58 3.01 6.86 ;
  LAYER M2 ;
        RECT 3.87 6.58 6.45 6.86 ;
  LAYER M2 ;
        RECT 7.31 6.58 8.17 6.86 ;
  LAYER M2 ;
        RECT 9.03 6.58 11.61 6.86 ;
  LAYER M2 ;
        RECT 12.47 6.58 13.33 6.86 ;
  LAYER M2 ;
        RECT 6.28 0.28 7.48 0.56 ;
  LAYER M2 ;
        RECT 11.01 0.7 12.21 0.98 ;
  LAYER M2 ;
        RECT 7.15 0.28 7.47 0.56 ;
  LAYER M1 ;
        RECT 7.185 0 7.435 0.42 ;
  LAYER M2 ;
        RECT 7.31 -0.14 10.75 0.14 ;
  LAYER M1 ;
        RECT 10.625 0 10.875 0.84 ;
  LAYER M2 ;
        RECT 10.75 0.7 11.18 0.98 ;
  LAYER M1 ;
        RECT 7.185 -0.085 7.435 0.085 ;
  LAYER M2 ;
        RECT 7.14 -0.14 7.48 0.14 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 0.505 ;
  LAYER M2 ;
        RECT 7.14 0.28 7.48 0.56 ;
  LAYER M1 ;
        RECT 10.625 -0.085 10.875 0.085 ;
  LAYER M2 ;
        RECT 10.58 -0.14 10.92 0.14 ;
  LAYER M1 ;
        RECT 10.625 0.755 10.875 0.925 ;
  LAYER M2 ;
        RECT 10.58 0.7 10.92 0.98 ;
  LAYER M1 ;
        RECT 7.185 -0.085 7.435 0.085 ;
  LAYER M2 ;
        RECT 7.14 -0.14 7.48 0.14 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 0.505 ;
  LAYER M2 ;
        RECT 7.14 0.28 7.48 0.56 ;
  LAYER M1 ;
        RECT 10.625 -0.085 10.875 0.085 ;
  LAYER M2 ;
        RECT 10.58 -0.14 10.92 0.14 ;
  LAYER M1 ;
        RECT 10.625 0.755 10.875 0.925 ;
  LAYER M2 ;
        RECT 10.58 0.7 10.92 0.98 ;
  LAYER M2 ;
        RECT 1.12 0.28 2.32 0.56 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M2 ;
        RECT 1.99 0.28 2.31 0.56 ;
  LAYER M1 ;
        RECT 2.025 0 2.275 0.42 ;
  LAYER M2 ;
        RECT 2.15 -0.14 5.59 0.14 ;
  LAYER M1 ;
        RECT 5.465 0 5.715 0.84 ;
  LAYER M2 ;
        RECT 5.59 0.7 6.02 0.98 ;
  LAYER M1 ;
        RECT 2.025 -0.085 2.275 0.085 ;
  LAYER M2 ;
        RECT 1.98 -0.14 2.32 0.14 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 0.505 ;
  LAYER M2 ;
        RECT 1.98 0.28 2.32 0.56 ;
  LAYER M1 ;
        RECT 5.465 -0.085 5.715 0.085 ;
  LAYER M2 ;
        RECT 5.42 -0.14 5.76 0.14 ;
  LAYER M1 ;
        RECT 5.465 0.755 5.715 0.925 ;
  LAYER M2 ;
        RECT 5.42 0.7 5.76 0.98 ;
  LAYER M1 ;
        RECT 2.025 -0.085 2.275 0.085 ;
  LAYER M2 ;
        RECT 1.98 -0.14 2.32 0.14 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 0.505 ;
  LAYER M2 ;
        RECT 1.98 0.28 2.32 0.56 ;
  LAYER M1 ;
        RECT 5.465 -0.085 5.715 0.085 ;
  LAYER M2 ;
        RECT 5.42 -0.14 5.76 0.14 ;
  LAYER M1 ;
        RECT 5.465 0.755 5.715 0.925 ;
  LAYER M2 ;
        RECT 5.42 0.7 5.76 0.98 ;
  LAYER M2 ;
        RECT 11.44 0.28 12.64 0.56 ;
  LAYER M2 ;
        RECT 13.59 0.7 14.79 0.98 ;
  LAYER M2 ;
        RECT 12.31 0.28 12.63 0.56 ;
  LAYER M1 ;
        RECT 12.345 0 12.595 0.42 ;
  LAYER M2 ;
        RECT 12.47 -0.14 13.33 0.14 ;
  LAYER M1 ;
        RECT 13.205 0 13.455 0.84 ;
  LAYER M2 ;
        RECT 13.33 0.7 13.76 0.98 ;
  LAYER M1 ;
        RECT 12.345 -0.085 12.595 0.085 ;
  LAYER M2 ;
        RECT 12.3 -0.14 12.64 0.14 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 0.505 ;
  LAYER M2 ;
        RECT 12.3 0.28 12.64 0.56 ;
  LAYER M1 ;
        RECT 13.205 -0.085 13.455 0.085 ;
  LAYER M2 ;
        RECT 13.16 -0.14 13.5 0.14 ;
  LAYER M1 ;
        RECT 13.205 0.755 13.455 0.925 ;
  LAYER M2 ;
        RECT 13.16 0.7 13.5 0.98 ;
  LAYER M1 ;
        RECT 12.345 -0.085 12.595 0.085 ;
  LAYER M2 ;
        RECT 12.3 -0.14 12.64 0.14 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 0.505 ;
  LAYER M2 ;
        RECT 12.3 0.28 12.64 0.56 ;
  LAYER M1 ;
        RECT 13.205 -0.085 13.455 0.085 ;
  LAYER M2 ;
        RECT 13.16 -0.14 13.5 0.14 ;
  LAYER M1 ;
        RECT 13.205 0.755 13.455 0.925 ;
  LAYER M2 ;
        RECT 13.16 0.7 13.5 0.98 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 8 0.28 9.2 0.56 ;
  LAYER M2 ;
        RECT 4.3 0.7 4.73 0.98 ;
  LAYER M1 ;
        RECT 4.605 0.84 4.855 1.26 ;
  LAYER M2 ;
        RECT 4.73 1.12 8.17 1.4 ;
  LAYER M1 ;
        RECT 8.045 0.42 8.295 1.26 ;
  LAYER M2 ;
        RECT 8.01 0.28 8.33 0.56 ;
  LAYER M1 ;
        RECT 4.605 0.755 4.855 0.925 ;
  LAYER M2 ;
        RECT 4.56 0.7 4.9 0.98 ;
  LAYER M1 ;
        RECT 4.605 1.175 4.855 1.345 ;
  LAYER M2 ;
        RECT 4.56 1.12 4.9 1.4 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 0.505 ;
  LAYER M2 ;
        RECT 8 0.28 8.34 0.56 ;
  LAYER M1 ;
        RECT 8.045 1.175 8.295 1.345 ;
  LAYER M2 ;
        RECT 8 1.12 8.34 1.4 ;
  LAYER M1 ;
        RECT 4.605 0.755 4.855 0.925 ;
  LAYER M2 ;
        RECT 4.56 0.7 4.9 0.98 ;
  LAYER M1 ;
        RECT 4.605 1.175 4.855 1.345 ;
  LAYER M2 ;
        RECT 4.56 1.12 4.9 1.4 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 0.505 ;
  LAYER M2 ;
        RECT 8 0.28 8.34 0.56 ;
  LAYER M1 ;
        RECT 8.045 1.175 8.295 1.345 ;
  LAYER M2 ;
        RECT 8 1.12 8.34 1.4 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M2 ;
        RECT 13.16 0.28 14.36 0.56 ;
  LAYER M2 ;
        RECT 9.46 0.7 9.89 0.98 ;
  LAYER M1 ;
        RECT 9.765 0.84 10.015 1.26 ;
  LAYER M2 ;
        RECT 9.89 1.12 13.33 1.4 ;
  LAYER M3 ;
        RECT 13.19 0.42 13.47 1.26 ;
  LAYER M2 ;
        RECT 13.17 0.28 13.49 0.56 ;
  LAYER M1 ;
        RECT 9.765 0.755 10.015 0.925 ;
  LAYER M2 ;
        RECT 9.72 0.7 10.06 0.98 ;
  LAYER M1 ;
        RECT 9.765 1.175 10.015 1.345 ;
  LAYER M2 ;
        RECT 9.72 1.12 10.06 1.4 ;
  LAYER M2 ;
        RECT 13.17 0.28 13.49 0.56 ;
  LAYER M3 ;
        RECT 13.19 0.26 13.47 0.58 ;
  LAYER M2 ;
        RECT 13.17 1.12 13.49 1.4 ;
  LAYER M3 ;
        RECT 13.19 1.1 13.47 1.42 ;
  LAYER M1 ;
        RECT 9.765 0.755 10.015 0.925 ;
  LAYER M2 ;
        RECT 9.72 0.7 10.06 0.98 ;
  LAYER M1 ;
        RECT 9.765 1.175 10.015 1.345 ;
  LAYER M2 ;
        RECT 9.72 1.12 10.06 1.4 ;
  LAYER M2 ;
        RECT 13.17 0.28 13.49 0.56 ;
  LAYER M3 ;
        RECT 13.19 0.26 13.47 0.58 ;
  LAYER M2 ;
        RECT 13.17 1.12 13.49 1.4 ;
  LAYER M3 ;
        RECT 13.19 1.1 13.47 1.42 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 2.84 0.28 4.04 0.56 ;
  LAYER M2 ;
        RECT 1.12 8.26 2.32 8.54 ;
  LAYER M2 ;
        RECT 2.84 8.26 4.04 8.54 ;
  LAYER M2 ;
        RECT 6.28 8.26 7.48 8.54 ;
  LAYER M2 ;
        RECT 8 8.26 9.2 8.54 ;
  LAYER M2 ;
        RECT 11.44 8.26 12.64 8.54 ;
  LAYER M2 ;
        RECT 13.16 8.26 14.36 8.54 ;
  LAYER M2 ;
        RECT 2.15 8.26 3.01 8.54 ;
  LAYER M2 ;
        RECT 3.87 8.26 6.45 8.54 ;
  LAYER M2 ;
        RECT 7.31 8.26 8.17 8.54 ;
  LAYER M2 ;
        RECT 9.03 8.26 11.61 8.54 ;
  LAYER M2 ;
        RECT 12.47 8.26 13.33 8.54 ;
  LAYER M2 ;
        RECT 11.44 14.56 12.64 14.84 ;
  LAYER M2 ;
        RECT 13.59 14.14 14.79 14.42 ;
  LAYER M2 ;
        RECT 12.31 14.56 12.63 14.84 ;
  LAYER M1 ;
        RECT 12.345 13.86 12.595 14.7 ;
  LAYER M2 ;
        RECT 12.47 13.72 13.33 14 ;
  LAYER M1 ;
        RECT 13.205 13.86 13.455 14.28 ;
  LAYER M2 ;
        RECT 13.33 14.14 13.76 14.42 ;
  LAYER M1 ;
        RECT 12.345 13.775 12.595 13.945 ;
  LAYER M2 ;
        RECT 12.3 13.72 12.64 14 ;
  LAYER M1 ;
        RECT 12.345 14.615 12.595 14.785 ;
  LAYER M2 ;
        RECT 12.3 14.56 12.64 14.84 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 13.945 ;
  LAYER M2 ;
        RECT 13.16 13.72 13.5 14 ;
  LAYER M1 ;
        RECT 13.205 14.195 13.455 14.365 ;
  LAYER M2 ;
        RECT 13.16 14.14 13.5 14.42 ;
  LAYER M1 ;
        RECT 12.345 13.775 12.595 13.945 ;
  LAYER M2 ;
        RECT 12.3 13.72 12.64 14 ;
  LAYER M1 ;
        RECT 12.345 14.615 12.595 14.785 ;
  LAYER M2 ;
        RECT 12.3 14.56 12.64 14.84 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 13.945 ;
  LAYER M2 ;
        RECT 13.16 13.72 13.5 14 ;
  LAYER M1 ;
        RECT 13.205 14.195 13.455 14.365 ;
  LAYER M2 ;
        RECT 13.16 14.14 13.5 14.42 ;
  LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
  LAYER M2 ;
        RECT 11.01 14.14 12.21 14.42 ;
  LAYER M2 ;
        RECT 7.15 14.56 7.47 14.84 ;
  LAYER M1 ;
        RECT 7.185 13.86 7.435 14.7 ;
  LAYER M2 ;
        RECT 7.31 13.72 10.75 14 ;
  LAYER M1 ;
        RECT 10.625 13.86 10.875 14.28 ;
  LAYER M2 ;
        RECT 10.75 14.14 11.18 14.42 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 13.945 ;
  LAYER M2 ;
        RECT 7.14 13.72 7.48 14 ;
  LAYER M1 ;
        RECT 7.185 14.615 7.435 14.785 ;
  LAYER M2 ;
        RECT 7.14 14.56 7.48 14.84 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 13.945 ;
  LAYER M2 ;
        RECT 10.58 13.72 10.92 14 ;
  LAYER M1 ;
        RECT 10.625 14.195 10.875 14.365 ;
  LAYER M2 ;
        RECT 10.58 14.14 10.92 14.42 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 13.945 ;
  LAYER M2 ;
        RECT 7.14 13.72 7.48 14 ;
  LAYER M1 ;
        RECT 7.185 14.615 7.435 14.785 ;
  LAYER M2 ;
        RECT 7.14 14.56 7.48 14.84 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 13.945 ;
  LAYER M2 ;
        RECT 10.58 13.72 10.92 14 ;
  LAYER M1 ;
        RECT 10.625 14.195 10.875 14.365 ;
  LAYER M2 ;
        RECT 10.58 14.14 10.92 14.42 ;
  LAYER M2 ;
        RECT 2.84 14.56 4.04 14.84 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 8 14.56 9.2 14.84 ;
  LAYER M2 ;
        RECT 4.3 14.14 5.16 14.42 ;
  LAYER M1 ;
        RECT 5.035 14.28 5.285 15.12 ;
  LAYER M2 ;
        RECT 5.16 14.98 8.17 15.26 ;
  LAYER M1 ;
        RECT 8.045 14.7 8.295 15.12 ;
  LAYER M2 ;
        RECT 8.01 14.56 8.33 14.84 ;
  LAYER M1 ;
        RECT 5.035 14.195 5.285 14.365 ;
  LAYER M2 ;
        RECT 4.99 14.14 5.33 14.42 ;
  LAYER M1 ;
        RECT 5.035 15.035 5.285 15.205 ;
  LAYER M2 ;
        RECT 4.99 14.98 5.33 15.26 ;
  LAYER M1 ;
        RECT 8.045 14.615 8.295 14.785 ;
  LAYER M2 ;
        RECT 8 14.56 8.34 14.84 ;
  LAYER M1 ;
        RECT 8.045 15.035 8.295 15.205 ;
  LAYER M2 ;
        RECT 8 14.98 8.34 15.26 ;
  LAYER M1 ;
        RECT 5.035 14.195 5.285 14.365 ;
  LAYER M2 ;
        RECT 4.99 14.14 5.33 14.42 ;
  LAYER M1 ;
        RECT 5.035 15.035 5.285 15.205 ;
  LAYER M2 ;
        RECT 4.99 14.98 5.33 15.26 ;
  LAYER M1 ;
        RECT 8.045 14.615 8.295 14.785 ;
  LAYER M2 ;
        RECT 8 14.56 8.34 14.84 ;
  LAYER M1 ;
        RECT 8.045 15.035 8.295 15.205 ;
  LAYER M2 ;
        RECT 8 14.98 8.34 15.26 ;
  LAYER M2 ;
        RECT 1.12 14.56 2.32 14.84 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 1.99 14.56 2.31 14.84 ;
  LAYER M1 ;
        RECT 2.025 13.86 2.275 14.7 ;
  LAYER M2 ;
        RECT 2.15 13.72 6.02 14 ;
  LAYER M3 ;
        RECT 5.88 13.86 6.16 14.28 ;
  LAYER M2 ;
        RECT 5.86 14.14 6.18 14.42 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 13.945 ;
  LAYER M2 ;
        RECT 1.98 13.72 2.32 14 ;
  LAYER M1 ;
        RECT 2.025 14.615 2.275 14.785 ;
  LAYER M2 ;
        RECT 1.98 14.56 2.32 14.84 ;
  LAYER M2 ;
        RECT 5.86 13.72 6.18 14 ;
  LAYER M3 ;
        RECT 5.88 13.7 6.16 14.02 ;
  LAYER M2 ;
        RECT 5.86 14.14 6.18 14.42 ;
  LAYER M3 ;
        RECT 5.88 14.12 6.16 14.44 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 13.945 ;
  LAYER M2 ;
        RECT 1.98 13.72 2.32 14 ;
  LAYER M1 ;
        RECT 2.025 14.615 2.275 14.785 ;
  LAYER M2 ;
        RECT 1.98 14.56 2.32 14.84 ;
  LAYER M2 ;
        RECT 5.86 13.72 6.18 14 ;
  LAYER M3 ;
        RECT 5.88 13.7 6.16 14.02 ;
  LAYER M2 ;
        RECT 5.86 14.14 6.18 14.42 ;
  LAYER M3 ;
        RECT 5.88 14.12 6.16 14.44 ;
  LAYER M2 ;
        RECT 8.43 14.14 9.63 14.42 ;
  LAYER M2 ;
        RECT 13.16 14.56 14.36 14.84 ;
  LAYER M2 ;
        RECT 9.46 14.14 9.89 14.42 ;
  LAYER M1 ;
        RECT 9.765 14.28 10.015 15.12 ;
  LAYER M2 ;
        RECT 9.89 14.98 13.33 15.26 ;
  LAYER M1 ;
        RECT 13.205 14.7 13.455 15.12 ;
  LAYER M2 ;
        RECT 13.17 14.56 13.49 14.84 ;
  LAYER M1 ;
        RECT 9.765 14.195 10.015 14.365 ;
  LAYER M2 ;
        RECT 9.72 14.14 10.06 14.42 ;
  LAYER M1 ;
        RECT 9.765 15.035 10.015 15.205 ;
  LAYER M2 ;
        RECT 9.72 14.98 10.06 15.26 ;
  LAYER M1 ;
        RECT 13.205 14.615 13.455 14.785 ;
  LAYER M2 ;
        RECT 13.16 14.56 13.5 14.84 ;
  LAYER M1 ;
        RECT 13.205 15.035 13.455 15.205 ;
  LAYER M2 ;
        RECT 13.16 14.98 13.5 15.26 ;
  LAYER M1 ;
        RECT 9.765 14.195 10.015 14.365 ;
  LAYER M2 ;
        RECT 9.72 14.14 10.06 14.42 ;
  LAYER M1 ;
        RECT 9.765 15.035 10.015 15.205 ;
  LAYER M2 ;
        RECT 9.72 14.98 10.06 15.26 ;
  LAYER M1 ;
        RECT 13.205 14.615 13.455 14.785 ;
  LAYER M2 ;
        RECT 13.16 14.56 13.5 14.84 ;
  LAYER M1 ;
        RECT 13.205 15.035 13.455 15.205 ;
  LAYER M2 ;
        RECT 13.16 14.98 13.5 15.26 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 3.865 ;
  LAYER M1 ;
        RECT 6.325 4.115 6.575 5.125 ;
  LAYER M1 ;
        RECT 6.325 6.215 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.755 0.335 7.005 3.865 ;
  LAYER M1 ;
        RECT 5.895 0.335 6.145 3.865 ;
  LAYER M2 ;
        RECT 6.28 6.58 7.48 6.86 ;
  LAYER M2 ;
        RECT 6.28 0.28 7.48 0.56 ;
  LAYER M2 ;
        RECT 6.28 4.48 7.48 4.76 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 3.865 ;
  LAYER M1 ;
        RECT 11.485 4.115 11.735 5.125 ;
  LAYER M1 ;
        RECT 11.485 6.215 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.915 0.335 12.165 3.865 ;
  LAYER M1 ;
        RECT 11.055 0.335 11.305 3.865 ;
  LAYER M2 ;
        RECT 11.44 6.58 12.64 6.86 ;
  LAYER M2 ;
        RECT 11.44 0.28 12.64 0.56 ;
  LAYER M2 ;
        RECT 11.44 4.48 12.64 4.76 ;
  LAYER M2 ;
        RECT 11.01 0.7 12.21 0.98 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 3.865 ;
  LAYER M1 ;
        RECT 8.905 4.115 9.155 5.125 ;
  LAYER M1 ;
        RECT 8.905 6.215 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.475 0.335 8.725 3.865 ;
  LAYER M1 ;
        RECT 9.335 0.335 9.585 3.865 ;
  LAYER M2 ;
        RECT 8 6.58 9.2 6.86 ;
  LAYER M2 ;
        RECT 8 0.28 9.2 0.56 ;
  LAYER M2 ;
        RECT 8 4.48 9.2 4.76 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 3.865 ;
  LAYER M1 ;
        RECT 14.065 4.115 14.315 5.125 ;
  LAYER M1 ;
        RECT 14.065 6.215 14.315 7.225 ;
  LAYER M1 ;
        RECT 13.635 0.335 13.885 3.865 ;
  LAYER M1 ;
        RECT 14.495 0.335 14.745 3.865 ;
  LAYER M2 ;
        RECT 13.16 6.58 14.36 6.86 ;
  LAYER M2 ;
        RECT 13.16 0.28 14.36 0.56 ;
  LAYER M2 ;
        RECT 13.16 4.48 14.36 4.76 ;
  LAYER M2 ;
        RECT 13.59 0.7 14.79 0.98 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 3.865 ;
  LAYER M1 ;
        RECT 1.165 4.115 1.415 5.125 ;
  LAYER M1 ;
        RECT 1.165 6.215 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.595 0.335 1.845 3.865 ;
  LAYER M1 ;
        RECT 0.735 0.335 0.985 3.865 ;
  LAYER M2 ;
        RECT 1.12 6.58 2.32 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.28 2.32 0.56 ;
  LAYER M2 ;
        RECT 1.12 4.48 2.32 4.76 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 3.865 ;
  LAYER M1 ;
        RECT 3.745 4.115 3.995 5.125 ;
  LAYER M1 ;
        RECT 3.745 6.215 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.315 0.335 3.565 3.865 ;
  LAYER M1 ;
        RECT 4.175 0.335 4.425 3.865 ;
  LAYER M2 ;
        RECT 2.84 6.58 4.04 6.86 ;
  LAYER M2 ;
        RECT 2.84 0.28 4.04 0.56 ;
  LAYER M2 ;
        RECT 2.84 4.48 4.04 4.76 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M1 ;
        RECT 11.485 11.255 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.485 9.995 11.735 11.005 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 8.905 ;
  LAYER M1 ;
        RECT 11.915 11.255 12.165 14.785 ;
  LAYER M1 ;
        RECT 11.055 11.255 11.305 14.785 ;
  LAYER M2 ;
        RECT 11.44 8.26 12.64 8.54 ;
  LAYER M2 ;
        RECT 11.44 14.56 12.64 14.84 ;
  LAYER M2 ;
        RECT 11.44 10.36 12.64 10.64 ;
  LAYER M2 ;
        RECT 11.01 14.14 12.21 14.42 ;
  LAYER M1 ;
        RECT 3.745 11.255 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.745 9.995 3.995 11.005 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 8.905 ;
  LAYER M1 ;
        RECT 3.315 11.255 3.565 14.785 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M2 ;
        RECT 2.84 8.26 4.04 8.54 ;
  LAYER M2 ;
        RECT 2.84 14.56 4.04 14.84 ;
  LAYER M2 ;
        RECT 2.84 10.36 4.04 10.64 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M2 ;
        RECT 6.28 8.26 7.48 8.54 ;
  LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
  LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M1 ;
        RECT 8.905 11.255 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.905 9.995 9.155 11.005 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 8.905 ;
  LAYER M1 ;
        RECT 8.475 11.255 8.725 14.785 ;
  LAYER M1 ;
        RECT 9.335 11.255 9.585 14.785 ;
  LAYER M2 ;
        RECT 8 8.26 9.2 8.54 ;
  LAYER M2 ;
        RECT 8 14.56 9.2 14.84 ;
  LAYER M2 ;
        RECT 8 10.36 9.2 10.64 ;
  LAYER M2 ;
        RECT 8.43 14.14 9.63 14.42 ;
  LAYER M1 ;
        RECT 14.065 11.255 14.315 14.785 ;
  LAYER M1 ;
        RECT 14.065 9.995 14.315 11.005 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 8.905 ;
  LAYER M1 ;
        RECT 13.635 11.255 13.885 14.785 ;
  LAYER M1 ;
        RECT 14.495 11.255 14.745 14.785 ;
  LAYER M2 ;
        RECT 13.16 8.26 14.36 8.54 ;
  LAYER M2 ;
        RECT 13.16 14.56 14.36 14.84 ;
  LAYER M2 ;
        RECT 13.16 10.36 14.36 10.64 ;
  LAYER M2 ;
        RECT 13.59 14.14 14.79 14.42 ;
  LAYER M1 ;
        RECT 1.165 11.255 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.165 9.995 1.415 11.005 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 8.905 ;
  LAYER M1 ;
        RECT 1.595 11.255 1.845 14.785 ;
  LAYER M1 ;
        RECT 0.735 11.255 0.985 14.785 ;
  LAYER M2 ;
        RECT 1.12 8.26 2.32 8.54 ;
  LAYER M2 ;
        RECT 1.12 14.56 2.32 14.84 ;
  LAYER M2 ;
        RECT 1.12 10.36 2.32 10.64 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  END 
END SECTION7
