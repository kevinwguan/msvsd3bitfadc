* NGSPICE file created from fn_postlayout.ext - technology: sky130A

*.subckt fn_postlayout a b c d e f vdd gnd
X0 a_44_18# c a_28_18# a_8_0# nmos
X1 a_60_76# e a_44_76# w_0_64# pmos
X2 a_44_76# c a_28_76# w_0_64# pmos
X3 a_92_18# d a_76_18# a_8_0# nmos
X4 a_76_18# f a_60_18# a_8_0# nmos
X5 a_28_18# a a_12_18# a_8_0# nmos
X6 a_108_18# b a_92_18# a_8_0# nmos
X7 a_92_76# d a_76_76# w_0_64# pmos
X8 a_76_76# f a_60_76# w_0_64# pmos
X9 a_28_76# a a_12_76# w_0_64# pmos
X10 a_108_76# b a_92_76# w_0_64# pmos
X11 a_60_18# e a_44_18# a_8_0# nmos
C0 a c 0.05fF
C1 b d 0.05fF
C2 f d 0.05fF
C3 e c 0.05fF
C4 f e 0.05fF
C5 m1_38_32# out 0.02fF
C6 out a_8_0# 0.01fF $ **FLOATING
C7 b a_8_0# 0.02fF
C8 a a_8_0# 0.02fF
C9 w_0_64# a_8_0# 0.05fF
*.ends

*X1 a b c d e f vdd gnd fn_postlayout
Vdd vdd gnd 2.5
V1 a gnd 0 pulse 0 2.5 0.1n 10p 10p 1n 2n
V2 b gnd 0 pulse 0 2.5 0.2n 10p 10p 1n 2n
V3 c gnd 0 pulse 0 2.5 0.3n 10p 10p 1n 2n
V4 d gnd 0 pulse 0 2.5 0.4n 10p 10p 1n 2n
V5 e gnd 0 pulse 0 2.5 0.5n 10p 10p 1n 2n
V6 f gnd 0 pulse 0 2.5 0.6n 10p 10p 1n 2n

***Simulation commands***
.op
.tran 10p 4n

*** .include model file ***
.include cmos.spice
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.end

