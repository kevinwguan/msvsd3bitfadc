MACRO STAGE2_INV_85542588
  ORIGIN 0 0 ;
  FOREIGN STAGE2_INV_85542588 0 0 ;
  SIZE 18.92 BY 21 ;
  PIN VI
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 15.34 2.78 15.62 8.98 ;
      LAYER M2 ;
        RECT 15.31 17.92 16.51 18.2 ;
      LAYER M3 ;
        RECT 15.34 8.82 15.62 18.06 ;
      LAYER M2 ;
        RECT 15.32 17.92 15.64 18.2 ;
    END
  END VI
  PIN SN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 14.12 6.59 20.32 ;
      LAYER M3 ;
        RECT 14.91 14.12 15.19 20.32 ;
      LAYER M3 ;
        RECT 6.31 14.515 6.59 14.885 ;
      LAYER M2 ;
        RECT 6.45 14.56 15.05 14.84 ;
      LAYER M3 ;
        RECT 14.91 14.515 15.19 14.885 ;
    END
  END SN
  PIN VO
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 5.45 6.98 5.73 13.18 ;
      LAYER M2 ;
        RECT 4.99 13.72 6.19 14 ;
      LAYER M3 ;
        RECT 5.45 13.02 5.73 13.86 ;
      LAYER M2 ;
        RECT 5.43 13.72 5.75 14 ;
    END
  END VO
  PIN SP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 0.68 6.59 12.76 ;
      LAYER M3 ;
        RECT 14.91 0.68 15.19 12.76 ;
      LAYER M3 ;
        RECT 6.31 1.075 6.59 1.445 ;
      LAYER M2 ;
        RECT 6.45 1.12 15.05 1.4 ;
      LAYER M3 ;
        RECT 14.91 1.075 15.19 1.445 ;
    END
  END SP
  OBS 
  LAYER M3 ;
        RECT 5.88 2.78 6.16 8.98 ;
  LAYER M2 ;
        RECT 4.99 17.92 6.19 18.2 ;
  LAYER M3 ;
        RECT 15.77 6.98 16.05 13.18 ;
  LAYER M2 ;
        RECT 15.31 13.72 16.51 14 ;
  LAYER M3 ;
        RECT 5.88 8.82 6.16 18.06 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 7.375 6.16 7.745 ;
  LAYER M2 ;
        RECT 6.02 7.42 15.91 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.375 16.05 7.745 ;
  LAYER M3 ;
        RECT 15.77 13.02 16.05 13.86 ;
  LAYER M2 ;
        RECT 15.75 13.72 16.07 14 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 15.75 7.42 16.07 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.4 16.05 7.72 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 15.75 7.42 16.07 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.4 16.05 7.72 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 15.75 7.42 16.07 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.4 16.05 7.72 ;
  LAYER M2 ;
        RECT 15.75 13.72 16.07 14 ;
  LAYER M3 ;
        RECT 15.77 13.7 16.05 14.02 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 15.75 7.42 16.07 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.4 16.05 7.72 ;
  LAYER M2 ;
        RECT 15.75 13.72 16.07 14 ;
  LAYER M3 ;
        RECT 15.77 13.7 16.05 14.02 ;
  LAYER M1 ;
        RECT 15.355 13.775 15.605 17.305 ;
  LAYER M1 ;
        RECT 15.355 17.555 15.605 18.565 ;
  LAYER M1 ;
        RECT 15.355 19.655 15.605 20.665 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 17.305 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 17.305 ;
  LAYER M2 ;
        RECT 14.88 14.14 16.08 14.42 ;
  LAYER M2 ;
        RECT 14.88 20.02 16.08 20.3 ;
  LAYER M2 ;
        RECT 15.31 13.72 16.51 14 ;
  LAYER M2 ;
        RECT 15.31 17.92 16.51 18.2 ;
  LAYER M3 ;
        RECT 14.91 14.12 15.19 20.32 ;
  LAYER M1 ;
        RECT 5.895 13.775 6.145 17.305 ;
  LAYER M1 ;
        RECT 5.895 17.555 6.145 18.565 ;
  LAYER M1 ;
        RECT 5.895 19.655 6.145 20.665 ;
  LAYER M1 ;
        RECT 5.465 13.775 5.715 17.305 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 17.305 ;
  LAYER M2 ;
        RECT 5.42 14.14 6.62 14.42 ;
  LAYER M2 ;
        RECT 5.42 20.02 6.62 20.3 ;
  LAYER M2 ;
        RECT 4.99 13.72 6.19 14 ;
  LAYER M2 ;
        RECT 4.99 17.92 6.19 18.2 ;
  LAYER M3 ;
        RECT 6.31 14.12 6.59 20.32 ;
  LAYER M1 ;
        RECT 17.505 9.575 17.755 13.105 ;
  LAYER M1 ;
        RECT 17.505 8.315 17.755 9.325 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 17.935 9.575 18.185 13.105 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M1 ;
        RECT 17.075 9.575 17.325 13.105 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.645 9.575 16.895 13.105 ;
  LAYER M1 ;
        RECT 16.645 8.315 16.895 9.325 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 16.215 9.575 16.465 13.105 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.785 9.575 16.035 13.105 ;
  LAYER M1 ;
        RECT 15.785 8.315 16.035 9.325 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 15.355 9.575 15.605 13.105 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 14.925 9.575 15.175 13.105 ;
  LAYER M1 ;
        RECT 14.925 8.315 15.175 9.325 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 9.575 14.745 13.105 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 14.065 9.575 14.315 13.105 ;
  LAYER M1 ;
        RECT 14.065 8.315 14.315 9.325 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 13.635 9.575 13.885 13.105 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 13.205 9.575 13.455 13.105 ;
  LAYER M1 ;
        RECT 13.205 8.315 13.455 9.325 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 9.575 13.025 13.105 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M2 ;
        RECT 13.16 12.88 17.8 13.16 ;
  LAYER M2 ;
        RECT 13.16 8.68 17.8 8.96 ;
  LAYER M2 ;
        RECT 12.73 12.46 18.23 12.74 ;
  LAYER M2 ;
        RECT 13.16 7 17.8 7.28 ;
  LAYER M2 ;
        RECT 13.16 2.8 17.8 3.08 ;
  LAYER M2 ;
        RECT 12.73 6.58 18.23 6.86 ;
  LAYER M2 ;
        RECT 13.16 0.7 17.8 0.98 ;
  LAYER M3 ;
        RECT 15.77 6.98 16.05 13.18 ;
  LAYER M3 ;
        RECT 15.34 2.78 15.62 8.98 ;
  LAYER M3 ;
        RECT 14.91 0.68 15.19 12.76 ;
  LAYER M1 ;
        RECT 1.165 9.575 1.415 13.105 ;
  LAYER M1 ;
        RECT 1.165 8.315 1.415 9.325 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 9.575 0.985 13.105 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 9.575 1.845 13.105 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 2.025 9.575 2.275 13.105 ;
  LAYER M1 ;
        RECT 2.025 8.315 2.275 9.325 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 9.575 2.705 13.105 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.885 9.575 3.135 13.105 ;
  LAYER M1 ;
        RECT 2.885 8.315 3.135 9.325 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 3.315 9.575 3.565 13.105 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 3.745 9.575 3.995 13.105 ;
  LAYER M1 ;
        RECT 3.745 8.315 3.995 9.325 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 9.575 4.425 13.105 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 4.605 9.575 4.855 13.105 ;
  LAYER M1 ;
        RECT 4.605 8.315 4.855 9.325 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 5.035 9.575 5.285 13.105 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.465 9.575 5.715 13.105 ;
  LAYER M1 ;
        RECT 5.465 8.315 5.715 9.325 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.895 9.575 6.145 13.105 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.325 9.575 6.575 13.105 ;
  LAYER M1 ;
        RECT 6.325 8.315 6.575 9.325 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 9.575 7.005 13.105 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 9.575 7.435 13.105 ;
  LAYER M1 ;
        RECT 7.185 8.315 7.435 9.325 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 9.575 7.865 13.105 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 8.045 9.575 8.295 13.105 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 9.325 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 8.475 9.575 8.725 13.105 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.905 9.575 9.155 13.105 ;
  LAYER M1 ;
        RECT 8.905 8.315 9.155 9.325 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 9.575 9.585 13.105 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 9.765 9.575 10.015 13.105 ;
  LAYER M1 ;
        RECT 9.765 8.315 10.015 9.325 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 10.195 9.575 10.445 13.105 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 10.625 9.575 10.875 13.105 ;
  LAYER M1 ;
        RECT 10.625 8.315 10.875 9.325 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 9.575 11.305 13.105 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M2 ;
        RECT 1.12 12.88 10.92 13.16 ;
  LAYER M2 ;
        RECT 1.12 8.68 10.92 8.96 ;
  LAYER M2 ;
        RECT 0.69 12.46 11.35 12.74 ;
  LAYER M2 ;
        RECT 1.12 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 10.92 3.08 ;
  LAYER M2 ;
        RECT 0.69 6.58 11.35 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.7 10.92 0.98 ;
  LAYER M3 ;
        RECT 5.45 6.98 5.73 13.18 ;
  LAYER M3 ;
        RECT 5.88 2.78 6.16 8.98 ;
  LAYER M3 ;
        RECT 6.31 0.68 6.59 12.76 ;
  END 
END STAGE2_INV_85542588
