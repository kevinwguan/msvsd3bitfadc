MACRO RING-FINAL
  ORIGIN 0 0 ;
  FOREIGN RING-FINAL 0 0 ;
  SIZE 57.62 BY 21 ;
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 14.12 6.59 20.32 ;
      LAYER M3 ;
        RECT 14.91 14.12 15.19 20.32 ;
      LAYER M3 ;
        RECT 6.31 14.515 6.59 14.885 ;
      LAYER M2 ;
        RECT 6.45 14.56 15.05 14.84 ;
      LAYER M3 ;
        RECT 14.91 14.515 15.19 14.885 ;
      LAYER M3 ;
        RECT 22.65 10.34 22.93 16.54 ;
      LAYER M3 ;
        RECT 27.38 10.34 27.66 16.54 ;
      LAYER M3 ;
        RECT 22.65 10.735 22.93 11.105 ;
      LAYER M2 ;
        RECT 22.79 10.78 27.52 11.06 ;
      LAYER M3 ;
        RECT 27.38 10.735 27.66 11.105 ;
      LAYER M2 ;
        RECT 31.22 10.78 32.42 11.06 ;
      LAYER M2 ;
        RECT 31.22 18.34 32.42 18.62 ;
      LAYER M3 ;
        RECT 34.26 14.12 34.54 20.32 ;
      LAYER M3 ;
        RECT 45.87 14.12 46.15 20.32 ;
      LAYER M2 ;
        RECT 15.05 14.56 22.79 14.84 ;
      LAYER M3 ;
        RECT 22.65 14.515 22.93 14.885 ;
      LAYER M2 ;
        RECT 27.52 10.78 31.39 11.06 ;
      LAYER M3 ;
        RECT 27.38 16.38 27.66 18.48 ;
      LAYER M2 ;
        RECT 27.52 18.34 31.39 18.62 ;
      LAYER M2 ;
        RECT 32.25 18.34 34.4 18.62 ;
      LAYER M3 ;
        RECT 34.26 18.295 34.54 18.665 ;
      LAYER M2 ;
        RECT 34.4 18.34 46.01 18.62 ;
      LAYER M3 ;
        RECT 45.87 18.295 46.15 18.665 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.31 0.68 6.59 12.76 ;
      LAYER M3 ;
        RECT 14.91 0.68 15.19 12.76 ;
      LAYER M3 ;
        RECT 6.31 1.075 6.59 1.445 ;
      LAYER M2 ;
        RECT 6.45 1.12 15.05 1.4 ;
      LAYER M3 ;
        RECT 14.91 1.075 15.19 1.445 ;
      LAYER M3 ;
        RECT 22.65 2.78 22.93 8.98 ;
      LAYER M3 ;
        RECT 27.38 2.78 27.66 8.98 ;
      LAYER M3 ;
        RECT 22.65 3.175 22.93 3.545 ;
      LAYER M2 ;
        RECT 22.79 3.22 27.52 3.5 ;
      LAYER M3 ;
        RECT 27.38 3.175 27.66 3.545 ;
      LAYER M2 ;
        RECT 31.22 4.48 32.42 4.76 ;
      LAYER M3 ;
        RECT 34.26 6.56 34.54 12.76 ;
      LAYER M3 ;
        RECT 45.87 0.68 46.15 12.76 ;
      LAYER M3 ;
        RECT 14.91 3.175 15.19 3.545 ;
      LAYER M2 ;
        RECT 15.05 3.22 22.79 3.5 ;
      LAYER M3 ;
        RECT 27.38 4.435 27.66 4.805 ;
      LAYER M2 ;
        RECT 27.52 4.48 31.39 4.76 ;
      LAYER M2 ;
        RECT 32.25 4.48 34.4 4.76 ;
      LAYER M3 ;
        RECT 34.26 4.62 34.54 6.72 ;
      LAYER M2 ;
        RECT 34.4 4.48 46.01 4.76 ;
      LAYER M3 ;
        RECT 45.87 4.435 46.15 4.805 ;
    END
  END VDD
  PIN CLKOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 31.22 12.04 32.42 12.32 ;
      LAYER M3 ;
        RECT 46.73 6.98 47.01 13.18 ;
      LAYER M2 ;
        RECT 46.27 13.72 47.47 14 ;
      LAYER M3 ;
        RECT 46.73 13.02 47.01 13.86 ;
      LAYER M2 ;
        RECT 46.71 13.72 47.03 14 ;
      LAYER M2 ;
        RECT 32.25 12.04 46.87 12.32 ;
      LAYER M3 ;
        RECT 46.73 11.995 47.01 12.365 ;
    END
  END CLKOUT
  PIN CLK1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 31.22 8.68 32.42 8.96 ;
      LAYER M2 ;
        RECT 32.94 8.68 34.14 8.96 ;
      LAYER M2 ;
        RECT 32.94 17.92 34.14 18.2 ;
      LAYER M2 ;
        RECT 32.95 8.68 33.27 8.96 ;
      LAYER M3 ;
        RECT 32.97 8.82 33.25 18.06 ;
      LAYER M2 ;
        RECT 32.95 17.92 33.27 18.2 ;
      LAYER M2 ;
        RECT 32.25 8.68 33.11 8.96 ;
    END
  END CLK1
  PIN CLK2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 32.94 12.88 34.14 13.16 ;
      LAYER M2 ;
        RECT 32.94 13.72 34.14 14 ;
      LAYER M2 ;
        RECT 32.95 12.88 33.27 13.16 ;
      LAYER M1 ;
        RECT 32.985 13.02 33.235 13.86 ;
      LAYER M2 ;
        RECT 32.95 13.72 33.27 14 ;
      LAYER M2 ;
        RECT 31.22 16.24 32.42 16.52 ;
      LAYER M1 ;
        RECT 32.985 13.86 33.235 16.38 ;
      LAYER M2 ;
        RECT 32.25 16.24 33.11 16.52 ;
    END
  END CLK2
  OBS 
  LAYER M2 ;
        RECT 26.92 4.9 28.98 5.18 ;
  LAYER M2 ;
        RECT 27.78 14.14 28.98 14.42 ;
  LAYER M2 ;
        RECT 28.22 4.9 28.54 5.18 ;
  LAYER M3 ;
        RECT 28.24 5.04 28.52 14.28 ;
  LAYER M2 ;
        RECT 28.22 14.14 28.54 14.42 ;
  LAYER M2 ;
        RECT 30.79 4.9 31.99 5.18 ;
  LAYER M2 ;
        RECT 30.79 12.46 31.99 12.74 ;
  LAYER M2 ;
        RECT 28.81 4.9 30.96 5.18 ;
  LAYER M3 ;
        RECT 28.24 12.415 28.52 12.785 ;
  LAYER M2 ;
        RECT 28.38 12.46 30.96 12.74 ;
  LAYER M2 ;
        RECT 28.22 12.46 28.54 12.74 ;
  LAYER M3 ;
        RECT 28.24 12.44 28.52 12.76 ;
  LAYER M2 ;
        RECT 28.22 12.46 28.54 12.74 ;
  LAYER M3 ;
        RECT 28.24 12.44 28.52 12.76 ;
  LAYER M3 ;
        RECT 15.34 2.78 15.62 8.98 ;
  LAYER M2 ;
        RECT 15.31 17.92 16.51 18.2 ;
  LAYER M3 ;
        RECT 15.34 8.82 15.62 18.06 ;
  LAYER M2 ;
        RECT 15.32 17.92 15.64 18.2 ;
  LAYER M2 ;
        RECT 20.04 9.1 24.68 9.38 ;
  LAYER M2 ;
        RECT 21.33 9.94 22.53 10.22 ;
  LAYER M2 ;
        RECT 21.77 9.1 22.09 9.38 ;
  LAYER M3 ;
        RECT 21.79 9.24 22.07 10.08 ;
  LAYER M2 ;
        RECT 21.77 9.94 22.09 10.22 ;
  LAYER M3 ;
        RECT 15.34 9.055 15.62 9.425 ;
  LAYER M2 ;
        RECT 15.48 9.1 20.21 9.38 ;
  LAYER M2 ;
        RECT 15.32 9.1 15.64 9.38 ;
  LAYER M3 ;
        RECT 15.34 9.08 15.62 9.4 ;
  LAYER M2 ;
        RECT 15.32 9.1 15.64 9.38 ;
  LAYER M3 ;
        RECT 15.34 9.08 15.62 9.4 ;
  LAYER M3 ;
        RECT 5.45 6.98 5.73 13.18 ;
  LAYER M2 ;
        RECT 4.99 13.72 6.19 14 ;
  LAYER M3 ;
        RECT 5.45 13.02 5.73 13.86 ;
  LAYER M2 ;
        RECT 5.43 13.72 5.75 14 ;
  LAYER M3 ;
        RECT 46.3 2.78 46.58 8.98 ;
  LAYER M2 ;
        RECT 46.27 17.92 47.47 18.2 ;
  LAYER M3 ;
        RECT 46.3 8.82 46.58 18.06 ;
  LAYER M2 ;
        RECT 46.28 17.92 46.6 18.2 ;
  LAYER M2 ;
        RECT 6.02 13.72 14.62 14 ;
  LAYER M3 ;
        RECT 14.48 13.739 14.76 13.981 ;
  LAYER M4 ;
        RECT 14.62 13.46 46.44 14.26 ;
  LAYER M3 ;
        RECT 46.3 13.675 46.58 14.045 ;
  LAYER M2 ;
        RECT 14.46 13.72 14.78 14 ;
  LAYER M3 ;
        RECT 14.48 13.7 14.76 14.02 ;
  LAYER M3 ;
        RECT 14.48 13.675 14.76 14.045 ;
  LAYER M4 ;
        RECT 14.455 13.46 14.785 14.26 ;
  LAYER M3 ;
        RECT 46.3 13.675 46.58 14.045 ;
  LAYER M4 ;
        RECT 46.275 13.46 46.605 14.26 ;
  LAYER M3 ;
        RECT 46.3 13.675 46.58 14.045 ;
  LAYER M4 ;
        RECT 46.275 13.46 46.605 14.26 ;
  LAYER M2 ;
        RECT 20.04 4.9 24.68 5.18 ;
  LAYER M2 ;
        RECT 21.33 14.14 22.53 14.42 ;
  LAYER M2 ;
        RECT 26.92 9.1 28.98 9.38 ;
  LAYER M2 ;
        RECT 27.78 9.94 28.98 10.22 ;
  LAYER M2 ;
        RECT 21.34 4.9 21.66 5.18 ;
  LAYER M3 ;
        RECT 21.36 5.04 21.64 14.28 ;
  LAYER M2 ;
        RECT 21.34 14.14 21.66 14.42 ;
  LAYER M3 ;
        RECT 21.36 9.475 21.64 9.845 ;
  LAYER M2 ;
        RECT 21.5 9.52 26.23 9.8 ;
  LAYER M1 ;
        RECT 26.105 9.24 26.355 9.66 ;
  LAYER M2 ;
        RECT 26.23 9.1 27.09 9.38 ;
  LAYER M2 ;
        RECT 27.79 9.1 28.11 9.38 ;
  LAYER M3 ;
        RECT 27.81 9.24 28.09 10.08 ;
  LAYER M2 ;
        RECT 27.79 9.94 28.11 10.22 ;
  LAYER M2 ;
        RECT 21.34 4.9 21.66 5.18 ;
  LAYER M3 ;
        RECT 21.36 4.88 21.64 5.2 ;
  LAYER M2 ;
        RECT 21.34 14.14 21.66 14.42 ;
  LAYER M3 ;
        RECT 21.36 14.12 21.64 14.44 ;
  LAYER M2 ;
        RECT 21.34 4.9 21.66 5.18 ;
  LAYER M3 ;
        RECT 21.36 4.88 21.64 5.2 ;
  LAYER M2 ;
        RECT 21.34 14.14 21.66 14.42 ;
  LAYER M3 ;
        RECT 21.36 14.12 21.64 14.44 ;
  LAYER M1 ;
        RECT 26.105 9.155 26.355 9.325 ;
  LAYER M2 ;
        RECT 26.06 9.1 26.4 9.38 ;
  LAYER M1 ;
        RECT 26.105 9.575 26.355 9.745 ;
  LAYER M2 ;
        RECT 26.06 9.52 26.4 9.8 ;
  LAYER M2 ;
        RECT 21.34 4.9 21.66 5.18 ;
  LAYER M3 ;
        RECT 21.36 4.88 21.64 5.2 ;
  LAYER M2 ;
        RECT 21.34 9.52 21.66 9.8 ;
  LAYER M3 ;
        RECT 21.36 9.5 21.64 9.82 ;
  LAYER M2 ;
        RECT 21.34 14.14 21.66 14.42 ;
  LAYER M3 ;
        RECT 21.36 14.12 21.64 14.44 ;
  LAYER M1 ;
        RECT 26.105 9.155 26.355 9.325 ;
  LAYER M2 ;
        RECT 26.06 9.1 26.4 9.38 ;
  LAYER M1 ;
        RECT 26.105 9.575 26.355 9.745 ;
  LAYER M2 ;
        RECT 26.06 9.52 26.4 9.8 ;
  LAYER M2 ;
        RECT 21.34 4.9 21.66 5.18 ;
  LAYER M3 ;
        RECT 21.36 4.88 21.64 5.2 ;
  LAYER M2 ;
        RECT 21.34 9.52 21.66 9.8 ;
  LAYER M3 ;
        RECT 21.36 9.5 21.64 9.82 ;
  LAYER M2 ;
        RECT 21.34 14.14 21.66 14.42 ;
  LAYER M3 ;
        RECT 21.36 14.12 21.64 14.44 ;
  LAYER M1 ;
        RECT 26.105 9.155 26.355 9.325 ;
  LAYER M2 ;
        RECT 26.06 9.1 26.4 9.38 ;
  LAYER M1 ;
        RECT 26.105 9.575 26.355 9.745 ;
  LAYER M2 ;
        RECT 26.06 9.52 26.4 9.8 ;
  LAYER M2 ;
        RECT 21.34 4.9 21.66 5.18 ;
  LAYER M3 ;
        RECT 21.36 4.88 21.64 5.2 ;
  LAYER M2 ;
        RECT 21.34 9.52 21.66 9.8 ;
  LAYER M3 ;
        RECT 21.36 9.5 21.64 9.82 ;
  LAYER M2 ;
        RECT 21.34 14.14 21.66 14.42 ;
  LAYER M3 ;
        RECT 21.36 14.12 21.64 14.44 ;
  LAYER M2 ;
        RECT 27.79 9.1 28.11 9.38 ;
  LAYER M3 ;
        RECT 27.81 9.08 28.09 9.4 ;
  LAYER M2 ;
        RECT 27.79 9.94 28.11 10.22 ;
  LAYER M3 ;
        RECT 27.81 9.92 28.09 10.24 ;
  LAYER M1 ;
        RECT 26.105 9.155 26.355 9.325 ;
  LAYER M2 ;
        RECT 26.06 9.1 26.4 9.38 ;
  LAYER M1 ;
        RECT 26.105 9.575 26.355 9.745 ;
  LAYER M2 ;
        RECT 26.06 9.52 26.4 9.8 ;
  LAYER M2 ;
        RECT 21.34 4.9 21.66 5.18 ;
  LAYER M3 ;
        RECT 21.36 4.88 21.64 5.2 ;
  LAYER M2 ;
        RECT 21.34 9.52 21.66 9.8 ;
  LAYER M3 ;
        RECT 21.36 9.5 21.64 9.82 ;
  LAYER M2 ;
        RECT 21.34 14.14 21.66 14.42 ;
  LAYER M3 ;
        RECT 21.36 14.12 21.64 14.44 ;
  LAYER M2 ;
        RECT 27.79 9.1 28.11 9.38 ;
  LAYER M3 ;
        RECT 27.81 9.08 28.09 9.4 ;
  LAYER M2 ;
        RECT 27.79 9.94 28.11 10.22 ;
  LAYER M3 ;
        RECT 27.81 9.92 28.09 10.24 ;
  LAYER M1 ;
        RECT 27.825 9.995 28.075 13.525 ;
  LAYER M1 ;
        RECT 27.825 13.775 28.075 14.785 ;
  LAYER M1 ;
        RECT 27.825 15.875 28.075 16.885 ;
  LAYER M1 ;
        RECT 28.255 9.995 28.505 13.525 ;
  LAYER M1 ;
        RECT 27.395 9.995 27.645 13.525 ;
  LAYER M2 ;
        RECT 27.35 10.36 28.55 10.64 ;
  LAYER M2 ;
        RECT 27.35 16.24 28.55 16.52 ;
  LAYER M2 ;
        RECT 27.78 9.94 28.98 10.22 ;
  LAYER M2 ;
        RECT 27.78 14.14 28.98 14.42 ;
  LAYER M3 ;
        RECT 27.38 10.34 27.66 16.54 ;
  LAYER M1 ;
        RECT 22.235 9.995 22.485 13.525 ;
  LAYER M1 ;
        RECT 22.235 13.775 22.485 14.785 ;
  LAYER M1 ;
        RECT 22.235 15.875 22.485 16.885 ;
  LAYER M1 ;
        RECT 21.805 9.995 22.055 13.525 ;
  LAYER M1 ;
        RECT 22.665 9.995 22.915 13.525 ;
  LAYER M2 ;
        RECT 21.76 10.36 22.96 10.64 ;
  LAYER M2 ;
        RECT 21.76 16.24 22.96 16.52 ;
  LAYER M2 ;
        RECT 21.33 9.94 22.53 10.22 ;
  LAYER M2 ;
        RECT 21.33 14.14 22.53 14.42 ;
  LAYER M3 ;
        RECT 22.65 10.34 22.93 16.54 ;
  LAYER M1 ;
        RECT 28.685 5.795 28.935 9.325 ;
  LAYER M1 ;
        RECT 28.685 4.535 28.935 5.545 ;
  LAYER M1 ;
        RECT 28.685 2.435 28.935 3.445 ;
  LAYER M1 ;
        RECT 29.115 5.795 29.365 9.325 ;
  LAYER M1 ;
        RECT 28.255 5.795 28.505 9.325 ;
  LAYER M1 ;
        RECT 27.825 5.795 28.075 9.325 ;
  LAYER M1 ;
        RECT 27.825 4.535 28.075 5.545 ;
  LAYER M1 ;
        RECT 27.825 2.435 28.075 3.445 ;
  LAYER M1 ;
        RECT 27.395 5.795 27.645 9.325 ;
  LAYER M1 ;
        RECT 26.965 5.795 27.215 9.325 ;
  LAYER M1 ;
        RECT 26.965 4.535 27.215 5.545 ;
  LAYER M1 ;
        RECT 26.965 2.435 27.215 3.445 ;
  LAYER M1 ;
        RECT 26.535 5.795 26.785 9.325 ;
  LAYER M2 ;
        RECT 26.49 8.68 29.41 8.96 ;
  LAYER M2 ;
        RECT 26.92 2.8 28.98 3.08 ;
  LAYER M2 ;
        RECT 26.92 9.1 28.98 9.38 ;
  LAYER M2 ;
        RECT 26.92 4.9 28.98 5.18 ;
  LAYER M3 ;
        RECT 27.38 2.78 27.66 8.98 ;
  LAYER M1 ;
        RECT 20.085 5.795 20.335 9.325 ;
  LAYER M1 ;
        RECT 20.085 4.535 20.335 5.545 ;
  LAYER M1 ;
        RECT 20.085 2.435 20.335 3.445 ;
  LAYER M1 ;
        RECT 19.655 5.795 19.905 9.325 ;
  LAYER M1 ;
        RECT 20.515 5.795 20.765 9.325 ;
  LAYER M1 ;
        RECT 20.945 5.795 21.195 9.325 ;
  LAYER M1 ;
        RECT 20.945 4.535 21.195 5.545 ;
  LAYER M1 ;
        RECT 20.945 2.435 21.195 3.445 ;
  LAYER M1 ;
        RECT 21.375 5.795 21.625 9.325 ;
  LAYER M1 ;
        RECT 21.805 5.795 22.055 9.325 ;
  LAYER M1 ;
        RECT 21.805 4.535 22.055 5.545 ;
  LAYER M1 ;
        RECT 21.805 2.435 22.055 3.445 ;
  LAYER M1 ;
        RECT 22.235 5.795 22.485 9.325 ;
  LAYER M1 ;
        RECT 22.665 5.795 22.915 9.325 ;
  LAYER M1 ;
        RECT 22.665 4.535 22.915 5.545 ;
  LAYER M1 ;
        RECT 22.665 2.435 22.915 3.445 ;
  LAYER M1 ;
        RECT 23.095 5.795 23.345 9.325 ;
  LAYER M1 ;
        RECT 23.525 5.795 23.775 9.325 ;
  LAYER M1 ;
        RECT 23.525 4.535 23.775 5.545 ;
  LAYER M1 ;
        RECT 23.525 2.435 23.775 3.445 ;
  LAYER M1 ;
        RECT 23.955 5.795 24.205 9.325 ;
  LAYER M1 ;
        RECT 24.385 5.795 24.635 9.325 ;
  LAYER M1 ;
        RECT 24.385 4.535 24.635 5.545 ;
  LAYER M1 ;
        RECT 24.385 2.435 24.635 3.445 ;
  LAYER M1 ;
        RECT 24.815 5.795 25.065 9.325 ;
  LAYER M2 ;
        RECT 19.61 8.68 25.11 8.96 ;
  LAYER M2 ;
        RECT 20.04 2.8 24.68 3.08 ;
  LAYER M2 ;
        RECT 20.04 9.1 24.68 9.38 ;
  LAYER M2 ;
        RECT 20.04 4.9 24.68 5.18 ;
  LAYER M3 ;
        RECT 22.65 2.78 22.93 8.98 ;
  LAYER M3 ;
        RECT 5.88 2.78 6.16 8.98 ;
  LAYER M2 ;
        RECT 4.99 17.92 6.19 18.2 ;
  LAYER M3 ;
        RECT 15.77 6.98 16.05 13.18 ;
  LAYER M2 ;
        RECT 15.31 13.72 16.51 14 ;
  LAYER M3 ;
        RECT 5.88 8.82 6.16 18.06 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 7.375 6.16 7.745 ;
  LAYER M2 ;
        RECT 6.02 7.42 15.91 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.375 16.05 7.745 ;
  LAYER M3 ;
        RECT 15.77 13.02 16.05 13.86 ;
  LAYER M2 ;
        RECT 15.75 13.72 16.07 14 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 15.75 7.42 16.07 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.4 16.05 7.72 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 15.75 7.42 16.07 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.4 16.05 7.72 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 15.75 7.42 16.07 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.4 16.05 7.72 ;
  LAYER M2 ;
        RECT 15.75 13.72 16.07 14 ;
  LAYER M3 ;
        RECT 15.77 13.7 16.05 14.02 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 17.92 6.18 18.2 ;
  LAYER M3 ;
        RECT 5.88 17.9 6.16 18.22 ;
  LAYER M2 ;
        RECT 15.75 7.42 16.07 7.7 ;
  LAYER M3 ;
        RECT 15.77 7.4 16.05 7.72 ;
  LAYER M2 ;
        RECT 15.75 13.72 16.07 14 ;
  LAYER M3 ;
        RECT 15.77 13.7 16.05 14.02 ;
  LAYER M1 ;
        RECT 15.355 13.775 15.605 17.305 ;
  LAYER M1 ;
        RECT 15.355 17.555 15.605 18.565 ;
  LAYER M1 ;
        RECT 15.355 19.655 15.605 20.665 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 17.305 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 17.305 ;
  LAYER M2 ;
        RECT 14.88 14.14 16.08 14.42 ;
  LAYER M2 ;
        RECT 14.88 20.02 16.08 20.3 ;
  LAYER M2 ;
        RECT 15.31 13.72 16.51 14 ;
  LAYER M2 ;
        RECT 15.31 17.92 16.51 18.2 ;
  LAYER M3 ;
        RECT 14.91 14.12 15.19 20.32 ;
  LAYER M1 ;
        RECT 5.895 13.775 6.145 17.305 ;
  LAYER M1 ;
        RECT 5.895 17.555 6.145 18.565 ;
  LAYER M1 ;
        RECT 5.895 19.655 6.145 20.665 ;
  LAYER M1 ;
        RECT 5.465 13.775 5.715 17.305 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 17.305 ;
  LAYER M2 ;
        RECT 5.42 14.14 6.62 14.42 ;
  LAYER M2 ;
        RECT 5.42 20.02 6.62 20.3 ;
  LAYER M2 ;
        RECT 4.99 13.72 6.19 14 ;
  LAYER M2 ;
        RECT 4.99 17.92 6.19 18.2 ;
  LAYER M3 ;
        RECT 6.31 14.12 6.59 20.32 ;
  LAYER M1 ;
        RECT 17.505 9.575 17.755 13.105 ;
  LAYER M1 ;
        RECT 17.505 8.315 17.755 9.325 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 17.935 9.575 18.185 13.105 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M1 ;
        RECT 17.075 9.575 17.325 13.105 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.645 9.575 16.895 13.105 ;
  LAYER M1 ;
        RECT 16.645 8.315 16.895 9.325 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 16.215 9.575 16.465 13.105 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.785 9.575 16.035 13.105 ;
  LAYER M1 ;
        RECT 15.785 8.315 16.035 9.325 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 15.355 9.575 15.605 13.105 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 14.925 9.575 15.175 13.105 ;
  LAYER M1 ;
        RECT 14.925 8.315 15.175 9.325 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 9.575 14.745 13.105 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 14.065 9.575 14.315 13.105 ;
  LAYER M1 ;
        RECT 14.065 8.315 14.315 9.325 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 13.635 9.575 13.885 13.105 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 13.205 9.575 13.455 13.105 ;
  LAYER M1 ;
        RECT 13.205 8.315 13.455 9.325 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 9.575 13.025 13.105 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M2 ;
        RECT 13.16 12.88 17.8 13.16 ;
  LAYER M2 ;
        RECT 13.16 8.68 17.8 8.96 ;
  LAYER M2 ;
        RECT 12.73 12.46 18.23 12.74 ;
  LAYER M2 ;
        RECT 13.16 7 17.8 7.28 ;
  LAYER M2 ;
        RECT 13.16 2.8 17.8 3.08 ;
  LAYER M2 ;
        RECT 12.73 6.58 18.23 6.86 ;
  LAYER M2 ;
        RECT 13.16 0.7 17.8 0.98 ;
  LAYER M3 ;
        RECT 15.77 6.98 16.05 13.18 ;
  LAYER M3 ;
        RECT 15.34 2.78 15.62 8.98 ;
  LAYER M3 ;
        RECT 14.91 0.68 15.19 12.76 ;
  LAYER M1 ;
        RECT 1.165 9.575 1.415 13.105 ;
  LAYER M1 ;
        RECT 1.165 8.315 1.415 9.325 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 9.575 0.985 13.105 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 9.575 1.845 13.105 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 2.025 9.575 2.275 13.105 ;
  LAYER M1 ;
        RECT 2.025 8.315 2.275 9.325 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 9.575 2.705 13.105 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.885 9.575 3.135 13.105 ;
  LAYER M1 ;
        RECT 2.885 8.315 3.135 9.325 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 3.315 9.575 3.565 13.105 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 3.745 9.575 3.995 13.105 ;
  LAYER M1 ;
        RECT 3.745 8.315 3.995 9.325 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 9.575 4.425 13.105 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 4.605 9.575 4.855 13.105 ;
  LAYER M1 ;
        RECT 4.605 8.315 4.855 9.325 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 5.035 9.575 5.285 13.105 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.465 9.575 5.715 13.105 ;
  LAYER M1 ;
        RECT 5.465 8.315 5.715 9.325 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.895 9.575 6.145 13.105 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.325 9.575 6.575 13.105 ;
  LAYER M1 ;
        RECT 6.325 8.315 6.575 9.325 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 9.575 7.005 13.105 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 9.575 7.435 13.105 ;
  LAYER M1 ;
        RECT 7.185 8.315 7.435 9.325 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 9.575 7.865 13.105 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 8.045 9.575 8.295 13.105 ;
  LAYER M1 ;
        RECT 8.045 8.315 8.295 9.325 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 8.475 9.575 8.725 13.105 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.905 9.575 9.155 13.105 ;
  LAYER M1 ;
        RECT 8.905 8.315 9.155 9.325 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 9.575 9.585 13.105 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 9.765 9.575 10.015 13.105 ;
  LAYER M1 ;
        RECT 9.765 8.315 10.015 9.325 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 10.195 9.575 10.445 13.105 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 10.625 9.575 10.875 13.105 ;
  LAYER M1 ;
        RECT 10.625 8.315 10.875 9.325 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 9.575 11.305 13.105 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M2 ;
        RECT 1.12 12.88 10.92 13.16 ;
  LAYER M2 ;
        RECT 1.12 8.68 10.92 8.96 ;
  LAYER M2 ;
        RECT 0.69 12.46 11.35 12.74 ;
  LAYER M2 ;
        RECT 1.12 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 10.92 3.08 ;
  LAYER M2 ;
        RECT 0.69 6.58 11.35 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.7 10.92 0.98 ;
  LAYER M3 ;
        RECT 5.45 6.98 5.73 13.18 ;
  LAYER M3 ;
        RECT 5.88 2.78 6.16 8.98 ;
  LAYER M3 ;
        RECT 6.31 0.68 6.59 12.76 ;
  LAYER M1 ;
        RECT 46.315 13.775 46.565 17.305 ;
  LAYER M1 ;
        RECT 46.315 17.555 46.565 18.565 ;
  LAYER M1 ;
        RECT 46.315 19.655 46.565 20.665 ;
  LAYER M1 ;
        RECT 46.745 13.775 46.995 17.305 ;
  LAYER M1 ;
        RECT 45.885 13.775 46.135 17.305 ;
  LAYER M2 ;
        RECT 45.84 14.14 47.04 14.42 ;
  LAYER M2 ;
        RECT 45.84 20.02 47.04 20.3 ;
  LAYER M2 ;
        RECT 46.27 13.72 47.47 14 ;
  LAYER M2 ;
        RECT 46.27 17.92 47.47 18.2 ;
  LAYER M3 ;
        RECT 45.87 14.12 46.15 20.32 ;
  LAYER M1 ;
        RECT 56.205 9.575 56.455 13.105 ;
  LAYER M1 ;
        RECT 56.205 8.315 56.455 9.325 ;
  LAYER M1 ;
        RECT 56.205 3.695 56.455 7.225 ;
  LAYER M1 ;
        RECT 56.205 2.435 56.455 3.445 ;
  LAYER M1 ;
        RECT 56.205 0.335 56.455 1.345 ;
  LAYER M1 ;
        RECT 56.635 9.575 56.885 13.105 ;
  LAYER M1 ;
        RECT 56.635 3.695 56.885 7.225 ;
  LAYER M1 ;
        RECT 55.775 9.575 56.025 13.105 ;
  LAYER M1 ;
        RECT 55.775 3.695 56.025 7.225 ;
  LAYER M1 ;
        RECT 55.345 9.575 55.595 13.105 ;
  LAYER M1 ;
        RECT 55.345 8.315 55.595 9.325 ;
  LAYER M1 ;
        RECT 55.345 3.695 55.595 7.225 ;
  LAYER M1 ;
        RECT 55.345 2.435 55.595 3.445 ;
  LAYER M1 ;
        RECT 55.345 0.335 55.595 1.345 ;
  LAYER M1 ;
        RECT 54.915 9.575 55.165 13.105 ;
  LAYER M1 ;
        RECT 54.915 3.695 55.165 7.225 ;
  LAYER M1 ;
        RECT 54.485 9.575 54.735 13.105 ;
  LAYER M1 ;
        RECT 54.485 8.315 54.735 9.325 ;
  LAYER M1 ;
        RECT 54.485 3.695 54.735 7.225 ;
  LAYER M1 ;
        RECT 54.485 2.435 54.735 3.445 ;
  LAYER M1 ;
        RECT 54.485 0.335 54.735 1.345 ;
  LAYER M1 ;
        RECT 54.055 9.575 54.305 13.105 ;
  LAYER M1 ;
        RECT 54.055 3.695 54.305 7.225 ;
  LAYER M1 ;
        RECT 53.625 9.575 53.875 13.105 ;
  LAYER M1 ;
        RECT 53.625 8.315 53.875 9.325 ;
  LAYER M1 ;
        RECT 53.625 3.695 53.875 7.225 ;
  LAYER M1 ;
        RECT 53.625 2.435 53.875 3.445 ;
  LAYER M1 ;
        RECT 53.625 0.335 53.875 1.345 ;
  LAYER M1 ;
        RECT 53.195 9.575 53.445 13.105 ;
  LAYER M1 ;
        RECT 53.195 3.695 53.445 7.225 ;
  LAYER M1 ;
        RECT 52.765 9.575 53.015 13.105 ;
  LAYER M1 ;
        RECT 52.765 8.315 53.015 9.325 ;
  LAYER M1 ;
        RECT 52.765 3.695 53.015 7.225 ;
  LAYER M1 ;
        RECT 52.765 2.435 53.015 3.445 ;
  LAYER M1 ;
        RECT 52.765 0.335 53.015 1.345 ;
  LAYER M1 ;
        RECT 52.335 9.575 52.585 13.105 ;
  LAYER M1 ;
        RECT 52.335 3.695 52.585 7.225 ;
  LAYER M1 ;
        RECT 51.905 9.575 52.155 13.105 ;
  LAYER M1 ;
        RECT 51.905 8.315 52.155 9.325 ;
  LAYER M1 ;
        RECT 51.905 3.695 52.155 7.225 ;
  LAYER M1 ;
        RECT 51.905 2.435 52.155 3.445 ;
  LAYER M1 ;
        RECT 51.905 0.335 52.155 1.345 ;
  LAYER M1 ;
        RECT 51.475 9.575 51.725 13.105 ;
  LAYER M1 ;
        RECT 51.475 3.695 51.725 7.225 ;
  LAYER M1 ;
        RECT 51.045 9.575 51.295 13.105 ;
  LAYER M1 ;
        RECT 51.045 8.315 51.295 9.325 ;
  LAYER M1 ;
        RECT 51.045 3.695 51.295 7.225 ;
  LAYER M1 ;
        RECT 51.045 2.435 51.295 3.445 ;
  LAYER M1 ;
        RECT 51.045 0.335 51.295 1.345 ;
  LAYER M1 ;
        RECT 50.615 9.575 50.865 13.105 ;
  LAYER M1 ;
        RECT 50.615 3.695 50.865 7.225 ;
  LAYER M1 ;
        RECT 50.185 9.575 50.435 13.105 ;
  LAYER M1 ;
        RECT 50.185 8.315 50.435 9.325 ;
  LAYER M1 ;
        RECT 50.185 3.695 50.435 7.225 ;
  LAYER M1 ;
        RECT 50.185 2.435 50.435 3.445 ;
  LAYER M1 ;
        RECT 50.185 0.335 50.435 1.345 ;
  LAYER M1 ;
        RECT 49.755 9.575 50.005 13.105 ;
  LAYER M1 ;
        RECT 49.755 3.695 50.005 7.225 ;
  LAYER M1 ;
        RECT 49.325 9.575 49.575 13.105 ;
  LAYER M1 ;
        RECT 49.325 8.315 49.575 9.325 ;
  LAYER M1 ;
        RECT 49.325 3.695 49.575 7.225 ;
  LAYER M1 ;
        RECT 49.325 2.435 49.575 3.445 ;
  LAYER M1 ;
        RECT 49.325 0.335 49.575 1.345 ;
  LAYER M1 ;
        RECT 48.895 9.575 49.145 13.105 ;
  LAYER M1 ;
        RECT 48.895 3.695 49.145 7.225 ;
  LAYER M1 ;
        RECT 48.465 9.575 48.715 13.105 ;
  LAYER M1 ;
        RECT 48.465 8.315 48.715 9.325 ;
  LAYER M1 ;
        RECT 48.465 3.695 48.715 7.225 ;
  LAYER M1 ;
        RECT 48.465 2.435 48.715 3.445 ;
  LAYER M1 ;
        RECT 48.465 0.335 48.715 1.345 ;
  LAYER M1 ;
        RECT 48.035 9.575 48.285 13.105 ;
  LAYER M1 ;
        RECT 48.035 3.695 48.285 7.225 ;
  LAYER M1 ;
        RECT 47.605 9.575 47.855 13.105 ;
  LAYER M1 ;
        RECT 47.605 8.315 47.855 9.325 ;
  LAYER M1 ;
        RECT 47.605 3.695 47.855 7.225 ;
  LAYER M1 ;
        RECT 47.605 2.435 47.855 3.445 ;
  LAYER M1 ;
        RECT 47.605 0.335 47.855 1.345 ;
  LAYER M1 ;
        RECT 47.175 9.575 47.425 13.105 ;
  LAYER M1 ;
        RECT 47.175 3.695 47.425 7.225 ;
  LAYER M1 ;
        RECT 46.745 9.575 46.995 13.105 ;
  LAYER M1 ;
        RECT 46.745 8.315 46.995 9.325 ;
  LAYER M1 ;
        RECT 46.745 3.695 46.995 7.225 ;
  LAYER M1 ;
        RECT 46.745 2.435 46.995 3.445 ;
  LAYER M1 ;
        RECT 46.745 0.335 46.995 1.345 ;
  LAYER M1 ;
        RECT 46.315 9.575 46.565 13.105 ;
  LAYER M1 ;
        RECT 46.315 3.695 46.565 7.225 ;
  LAYER M1 ;
        RECT 45.885 9.575 46.135 13.105 ;
  LAYER M1 ;
        RECT 45.885 8.315 46.135 9.325 ;
  LAYER M1 ;
        RECT 45.885 3.695 46.135 7.225 ;
  LAYER M1 ;
        RECT 45.885 2.435 46.135 3.445 ;
  LAYER M1 ;
        RECT 45.885 0.335 46.135 1.345 ;
  LAYER M1 ;
        RECT 45.455 9.575 45.705 13.105 ;
  LAYER M1 ;
        RECT 45.455 3.695 45.705 7.225 ;
  LAYER M1 ;
        RECT 45.025 9.575 45.275 13.105 ;
  LAYER M1 ;
        RECT 45.025 8.315 45.275 9.325 ;
  LAYER M1 ;
        RECT 45.025 3.695 45.275 7.225 ;
  LAYER M1 ;
        RECT 45.025 2.435 45.275 3.445 ;
  LAYER M1 ;
        RECT 45.025 0.335 45.275 1.345 ;
  LAYER M1 ;
        RECT 44.595 9.575 44.845 13.105 ;
  LAYER M1 ;
        RECT 44.595 3.695 44.845 7.225 ;
  LAYER M1 ;
        RECT 44.165 9.575 44.415 13.105 ;
  LAYER M1 ;
        RECT 44.165 8.315 44.415 9.325 ;
  LAYER M1 ;
        RECT 44.165 3.695 44.415 7.225 ;
  LAYER M1 ;
        RECT 44.165 2.435 44.415 3.445 ;
  LAYER M1 ;
        RECT 44.165 0.335 44.415 1.345 ;
  LAYER M1 ;
        RECT 43.735 9.575 43.985 13.105 ;
  LAYER M1 ;
        RECT 43.735 3.695 43.985 7.225 ;
  LAYER M1 ;
        RECT 43.305 9.575 43.555 13.105 ;
  LAYER M1 ;
        RECT 43.305 8.315 43.555 9.325 ;
  LAYER M1 ;
        RECT 43.305 3.695 43.555 7.225 ;
  LAYER M1 ;
        RECT 43.305 2.435 43.555 3.445 ;
  LAYER M1 ;
        RECT 43.305 0.335 43.555 1.345 ;
  LAYER M1 ;
        RECT 42.875 9.575 43.125 13.105 ;
  LAYER M1 ;
        RECT 42.875 3.695 43.125 7.225 ;
  LAYER M1 ;
        RECT 42.445 9.575 42.695 13.105 ;
  LAYER M1 ;
        RECT 42.445 8.315 42.695 9.325 ;
  LAYER M1 ;
        RECT 42.445 3.695 42.695 7.225 ;
  LAYER M1 ;
        RECT 42.445 2.435 42.695 3.445 ;
  LAYER M1 ;
        RECT 42.445 0.335 42.695 1.345 ;
  LAYER M1 ;
        RECT 42.015 9.575 42.265 13.105 ;
  LAYER M1 ;
        RECT 42.015 3.695 42.265 7.225 ;
  LAYER M1 ;
        RECT 41.585 9.575 41.835 13.105 ;
  LAYER M1 ;
        RECT 41.585 8.315 41.835 9.325 ;
  LAYER M1 ;
        RECT 41.585 3.695 41.835 7.225 ;
  LAYER M1 ;
        RECT 41.585 2.435 41.835 3.445 ;
  LAYER M1 ;
        RECT 41.585 0.335 41.835 1.345 ;
  LAYER M1 ;
        RECT 41.155 9.575 41.405 13.105 ;
  LAYER M1 ;
        RECT 41.155 3.695 41.405 7.225 ;
  LAYER M1 ;
        RECT 40.725 9.575 40.975 13.105 ;
  LAYER M1 ;
        RECT 40.725 8.315 40.975 9.325 ;
  LAYER M1 ;
        RECT 40.725 3.695 40.975 7.225 ;
  LAYER M1 ;
        RECT 40.725 2.435 40.975 3.445 ;
  LAYER M1 ;
        RECT 40.725 0.335 40.975 1.345 ;
  LAYER M1 ;
        RECT 40.295 9.575 40.545 13.105 ;
  LAYER M1 ;
        RECT 40.295 3.695 40.545 7.225 ;
  LAYER M1 ;
        RECT 39.865 9.575 40.115 13.105 ;
  LAYER M1 ;
        RECT 39.865 8.315 40.115 9.325 ;
  LAYER M1 ;
        RECT 39.865 3.695 40.115 7.225 ;
  LAYER M1 ;
        RECT 39.865 2.435 40.115 3.445 ;
  LAYER M1 ;
        RECT 39.865 0.335 40.115 1.345 ;
  LAYER M1 ;
        RECT 39.435 9.575 39.685 13.105 ;
  LAYER M1 ;
        RECT 39.435 3.695 39.685 7.225 ;
  LAYER M1 ;
        RECT 39.005 9.575 39.255 13.105 ;
  LAYER M1 ;
        RECT 39.005 8.315 39.255 9.325 ;
  LAYER M1 ;
        RECT 39.005 3.695 39.255 7.225 ;
  LAYER M1 ;
        RECT 39.005 2.435 39.255 3.445 ;
  LAYER M1 ;
        RECT 39.005 0.335 39.255 1.345 ;
  LAYER M1 ;
        RECT 38.575 9.575 38.825 13.105 ;
  LAYER M1 ;
        RECT 38.575 3.695 38.825 7.225 ;
  LAYER M1 ;
        RECT 38.145 9.575 38.395 13.105 ;
  LAYER M1 ;
        RECT 38.145 8.315 38.395 9.325 ;
  LAYER M1 ;
        RECT 38.145 3.695 38.395 7.225 ;
  LAYER M1 ;
        RECT 38.145 2.435 38.395 3.445 ;
  LAYER M1 ;
        RECT 38.145 0.335 38.395 1.345 ;
  LAYER M1 ;
        RECT 37.715 9.575 37.965 13.105 ;
  LAYER M1 ;
        RECT 37.715 3.695 37.965 7.225 ;
  LAYER M1 ;
        RECT 37.285 9.575 37.535 13.105 ;
  LAYER M1 ;
        RECT 37.285 8.315 37.535 9.325 ;
  LAYER M1 ;
        RECT 37.285 3.695 37.535 7.225 ;
  LAYER M1 ;
        RECT 37.285 2.435 37.535 3.445 ;
  LAYER M1 ;
        RECT 37.285 0.335 37.535 1.345 ;
  LAYER M1 ;
        RECT 36.855 9.575 37.105 13.105 ;
  LAYER M1 ;
        RECT 36.855 3.695 37.105 7.225 ;
  LAYER M1 ;
        RECT 36.425 9.575 36.675 13.105 ;
  LAYER M1 ;
        RECT 36.425 8.315 36.675 9.325 ;
  LAYER M1 ;
        RECT 36.425 3.695 36.675 7.225 ;
  LAYER M1 ;
        RECT 36.425 2.435 36.675 3.445 ;
  LAYER M1 ;
        RECT 36.425 0.335 36.675 1.345 ;
  LAYER M1 ;
        RECT 35.995 9.575 36.245 13.105 ;
  LAYER M1 ;
        RECT 35.995 3.695 36.245 7.225 ;
  LAYER M2 ;
        RECT 36.38 12.88 56.5 13.16 ;
  LAYER M2 ;
        RECT 36.38 8.68 56.5 8.96 ;
  LAYER M2 ;
        RECT 35.95 12.46 56.93 12.74 ;
  LAYER M2 ;
        RECT 36.38 7 56.5 7.28 ;
  LAYER M2 ;
        RECT 36.38 2.8 56.5 3.08 ;
  LAYER M2 ;
        RECT 35.95 6.58 56.93 6.86 ;
  LAYER M2 ;
        RECT 36.38 0.7 56.5 0.98 ;
  LAYER M3 ;
        RECT 46.73 6.98 47.01 13.18 ;
  LAYER M3 ;
        RECT 46.3 2.78 46.58 8.98 ;
  LAYER M3 ;
        RECT 45.87 0.68 46.15 12.76 ;
  LAYER M1 ;
        RECT 33.845 13.775 34.095 17.305 ;
  LAYER M1 ;
        RECT 33.845 17.555 34.095 18.565 ;
  LAYER M1 ;
        RECT 33.845 19.655 34.095 20.665 ;
  LAYER M1 ;
        RECT 33.415 13.775 33.665 17.305 ;
  LAYER M1 ;
        RECT 34.275 13.775 34.525 17.305 ;
  LAYER M2 ;
        RECT 33.37 14.14 34.57 14.42 ;
  LAYER M2 ;
        RECT 33.37 20.02 34.57 20.3 ;
  LAYER M2 ;
        RECT 32.94 13.72 34.14 14 ;
  LAYER M2 ;
        RECT 32.94 17.92 34.14 18.2 ;
  LAYER M3 ;
        RECT 34.26 14.12 34.54 20.32 ;
  LAYER M1 ;
        RECT 33.845 9.575 34.095 13.105 ;
  LAYER M1 ;
        RECT 33.845 8.315 34.095 9.325 ;
  LAYER M1 ;
        RECT 33.845 6.215 34.095 7.225 ;
  LAYER M1 ;
        RECT 33.415 9.575 33.665 13.105 ;
  LAYER M1 ;
        RECT 34.275 9.575 34.525 13.105 ;
  LAYER M2 ;
        RECT 33.37 12.46 34.57 12.74 ;
  LAYER M2 ;
        RECT 33.37 6.58 34.57 6.86 ;
  LAYER M2 ;
        RECT 32.94 12.88 34.14 13.16 ;
  LAYER M2 ;
        RECT 32.94 8.68 34.14 8.96 ;
  LAYER M3 ;
        RECT 34.26 6.56 34.54 12.76 ;
  LAYER M1 ;
        RECT 31.265 12.095 31.515 15.625 ;
  LAYER M1 ;
        RECT 31.265 15.875 31.515 16.885 ;
  LAYER M1 ;
        RECT 31.265 17.975 31.515 18.985 ;
  LAYER M1 ;
        RECT 31.695 12.095 31.945 15.625 ;
  LAYER M1 ;
        RECT 30.835 12.095 31.085 15.625 ;
  LAYER M2 ;
        RECT 31.22 18.34 32.42 18.62 ;
  LAYER M2 ;
        RECT 31.22 12.04 32.42 12.32 ;
  LAYER M2 ;
        RECT 31.22 16.24 32.42 16.52 ;
  LAYER M2 ;
        RECT 30.79 12.46 31.99 12.74 ;
  LAYER M1 ;
        RECT 31.265 4.535 31.515 8.065 ;
  LAYER M1 ;
        RECT 31.265 8.315 31.515 9.325 ;
  LAYER M1 ;
        RECT 31.265 10.415 31.515 11.425 ;
  LAYER M1 ;
        RECT 31.695 4.535 31.945 8.065 ;
  LAYER M1 ;
        RECT 30.835 4.535 31.085 8.065 ;
  LAYER M2 ;
        RECT 31.22 10.78 32.42 11.06 ;
  LAYER M2 ;
        RECT 31.22 4.48 32.42 4.76 ;
  LAYER M2 ;
        RECT 31.22 8.68 32.42 8.96 ;
  LAYER M2 ;
        RECT 30.79 4.9 31.99 5.18 ;
  END 
END RING-FINAL
