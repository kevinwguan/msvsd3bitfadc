MACRO COUNTER
  ORIGIN 0 0 ;
  FOREIGN COUNTER 0 0 ;
  SIZE 12.9 BY 15.12 ;
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
      LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
      LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
      LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
      LAYER M3 ;
        RECT 4.16 8.635 4.44 9.005 ;
      LAYER M2 ;
        RECT 4.3 8.68 6.02 8.96 ;
      LAYER M3 ;
        RECT 5.88 8.635 6.16 9.005 ;
      LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
      LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
      LAYER M3 ;
        RECT 11.04 0.68 11.32 6.88 ;
      LAYER M3 ;
        RECT 1.58 6.72 1.86 8.4 ;
      LAYER M3 ;
        RECT 1.58 8.635 1.86 9.005 ;
      LAYER M2 ;
        RECT 1.72 8.68 4.3 8.96 ;
      LAYER M2 ;
        RECT 6.02 8.68 9.46 8.96 ;
      LAYER M3 ;
        RECT 9.32 8.635 9.6 9.005 ;
      LAYER M2 ;
        RECT 9.46 8.68 11.18 8.96 ;
      LAYER M3 ;
        RECT 11.04 8.635 11.32 9.005 ;
      LAYER M3 ;
        RECT 11.04 6.72 11.32 8.4 ;
    END
  END GND
  PIN IN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
      LAYER M3 ;
        RECT 5.88 0.68 6.16 6.88 ;
      LAYER M3 ;
        RECT 4.16 1.075 4.44 1.445 ;
      LAYER M2 ;
        RECT 4.3 1.12 6.02 1.4 ;
      LAYER M3 ;
        RECT 5.88 1.075 6.16 1.445 ;
      LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
      LAYER M2 ;
        RECT 6.02 1.12 9.46 1.4 ;
      LAYER M3 ;
        RECT 9.32 1.075 9.6 1.445 ;
    END
  END IN
  PIN CLK
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 2.84 2.8 4.04 3.08 ;
      LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
      LAYER M2 ;
        RECT 2.85 2.8 3.17 3.08 ;
      LAYER M3 ;
        RECT 2.87 2.94 3.15 12.18 ;
      LAYER M2 ;
        RECT 2.85 12.04 3.17 12.32 ;
      LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
      LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
      LAYER M2 ;
        RECT 8.01 7 8.33 7.28 ;
      LAYER M1 ;
        RECT 8.045 7.14 8.295 7.98 ;
      LAYER M2 ;
        RECT 8.01 7.84 8.33 8.12 ;
      LAYER M3 ;
        RECT 2.87 7.375 3.15 7.745 ;
      LAYER M2 ;
        RECT 3.01 7.42 8.17 7.7 ;
      LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
    END
  END CLK
  PIN Q0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.15 7.82 1.43 12.34 ;
    END
  END Q0
  PIN Q3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.15 0.26 1.43 4.78 ;
    END
  END Q3
  PIN Q2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 11.47 0.26 11.75 4.78 ;
    END
  END Q2
  PIN Q1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 11.47 7.82 11.75 12.34 ;
    END
  END Q1
  OBS 
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M2 ;
        RECT 8.01 2.8 8.33 3.08 ;
  LAYER M3 ;
        RECT 8.03 2.94 8.31 12.18 ;
  LAYER M2 ;
        RECT 8.01 12.04 8.33 12.32 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M1 ;
        RECT 7.185 7.14 7.435 7.98 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 8.03 7.375 8.31 7.745 ;
  LAYER M4 ;
        RECT 7.31 7.16 8.17 7.96 ;
  LAYER M3 ;
        RECT 7.17 7.14 7.45 7.56 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 6.98 7.45 7.3 ;
  LAYER M3 ;
        RECT 7.17 7.375 7.45 7.745 ;
  LAYER M4 ;
        RECT 7.145 7.16 7.475 7.96 ;
  LAYER M3 ;
        RECT 8.03 7.375 8.31 7.745 ;
  LAYER M4 ;
        RECT 8.005 7.16 8.335 7.96 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 6.98 7.45 7.3 ;
  LAYER M3 ;
        RECT 7.17 7.375 7.45 7.745 ;
  LAYER M4 ;
        RECT 7.145 7.16 7.475 7.96 ;
  LAYER M3 ;
        RECT 8.03 7.375 8.31 7.745 ;
  LAYER M4 ;
        RECT 8.005 7.16 8.335 7.96 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 2.84 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M2 ;
        RECT 4.73 2.8 6.45 3.08 ;
  LAYER M1 ;
        RECT 4.605 2.94 4.855 7.14 ;
  LAYER M2 ;
        RECT 3.87 7 4.73 7.28 ;
  LAYER M2 ;
        RECT 2.85 7 3.17 7.28 ;
  LAYER M1 ;
        RECT 2.885 7.14 3.135 7.98 ;
  LAYER M2 ;
        RECT 2.85 7.84 3.17 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.14 4.855 12.18 ;
  LAYER M2 ;
        RECT 4.73 12.04 6.45 12.32 ;
  LAYER M1 ;
        RECT 4.605 2.855 4.855 3.025 ;
  LAYER M2 ;
        RECT 4.56 2.8 4.9 3.08 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 4.605 2.855 4.855 3.025 ;
  LAYER M2 ;
        RECT 4.56 2.8 4.9 3.08 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 2.885 7.055 3.135 7.225 ;
  LAYER M2 ;
        RECT 2.84 7 3.18 7.28 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 4.605 2.855 4.855 3.025 ;
  LAYER M2 ;
        RECT 4.56 2.8 4.9 3.08 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 2.885 7.055 3.135 7.225 ;
  LAYER M2 ;
        RECT 2.84 7 3.18 7.28 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 4.605 2.855 4.855 3.025 ;
  LAYER M2 ;
        RECT 4.56 2.8 4.9 3.08 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 2.885 7.055 3.135 7.225 ;
  LAYER M2 ;
        RECT 2.84 7 3.18 7.28 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 4.605 2.855 4.855 3.025 ;
  LAYER M2 ;
        RECT 4.56 2.8 4.9 3.08 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 4.605 12.095 4.855 12.265 ;
  LAYER M2 ;
        RECT 4.56 12.04 4.9 12.32 ;
  LAYER M1 ;
        RECT 2.885 7.055 3.135 7.225 ;
  LAYER M2 ;
        RECT 2.84 7 3.18 7.28 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 8.065 ;
  LAYER M2 ;
        RECT 2.84 7.84 3.18 8.12 ;
  LAYER M1 ;
        RECT 4.605 2.855 4.855 3.025 ;
  LAYER M2 ;
        RECT 4.56 2.8 4.9 3.08 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 4.605 12.095 4.855 12.265 ;
  LAYER M2 ;
        RECT 4.56 12.04 4.9 12.32 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 2.84 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 2.84 2.8 4.04 3.08 ;
  LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M2 ;
        RECT 5.85 6.58 7.05 6.86 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 6.88 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
  LAYER M2 ;
        RECT 8.43 14.14 9.63 14.42 ;
  LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 8.43 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M3 ;
        RECT 1.15 7.82 1.43 12.34 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 3.865 ;
  LAYER M1 ;
        RECT 1.165 4.115 1.415 5.125 ;
  LAYER M1 ;
        RECT 1.165 6.215 1.415 7.225 ;
  LAYER M1 ;
        RECT 0.735 0.335 0.985 3.865 ;
  LAYER M1 ;
        RECT 1.595 0.335 1.845 3.865 ;
  LAYER M2 ;
        RECT 0.26 0.28 1.46 0.56 ;
  LAYER M2 ;
        RECT 0.26 4.48 1.46 4.76 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M3 ;
        RECT 1.15 0.26 1.43 4.78 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 3.865 ;
  LAYER M1 ;
        RECT 11.485 4.115 11.735 5.125 ;
  LAYER M1 ;
        RECT 11.485 6.215 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.915 0.335 12.165 3.865 ;
  LAYER M1 ;
        RECT 11.055 0.335 11.305 3.865 ;
  LAYER M2 ;
        RECT 11.44 0.28 12.64 0.56 ;
  LAYER M2 ;
        RECT 11.44 4.48 12.64 4.76 ;
  LAYER M2 ;
        RECT 11.01 0.7 12.21 0.98 ;
  LAYER M2 ;
        RECT 11.01 6.58 12.21 6.86 ;
  LAYER M3 ;
        RECT 11.47 0.26 11.75 4.78 ;
  LAYER M3 ;
        RECT 11.04 0.68 11.32 6.88 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M2 ;
        RECT 11.44 7.84 12.64 8.12 ;
  LAYER M2 ;
        RECT 11.44 12.04 12.64 12.32 ;
  LAYER M2 ;
        RECT 11.01 8.26 12.21 8.54 ;
  LAYER M2 ;
        RECT 11.01 14.14 12.21 14.42 ;
  LAYER M3 ;
        RECT 11.47 7.82 11.75 12.34 ;
  LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
  END 
END COUNTER
