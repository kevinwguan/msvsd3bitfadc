MACRO PMOS_S_81354572_X2_Y3
  UNITS 
    DATABASE MICRONS UNITS 1000;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN PMOS_S_81354572_X2_Y3 0 0 ;
  SIZE 3440 BY 19320 ;
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1150 260 1430 12340 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1580 4460 1860 16540 ;
    END
  END G
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2010 680 2290 18640 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1165 335 1415 3865 ;
    LAYER M1 ;
      RECT 1165 4115 1415 5125 ;
    LAYER M1 ;
      RECT 1165 6215 1415 9745 ;
    LAYER M1 ;
      RECT 1165 9995 1415 11005 ;
    LAYER M1 ;
      RECT 1165 12095 1415 15625 ;
    LAYER M1 ;
      RECT 1165 15875 1415 16885 ;
    LAYER M1 ;
      RECT 1165 17975 1415 18985 ;
    LAYER M1 ;
      RECT 735 335 985 3865 ;
    LAYER M1 ;
      RECT 735 6215 985 9745 ;
    LAYER M1 ;
      RECT 735 12095 985 15625 ;
    LAYER M1 ;
      RECT 1595 335 1845 3865 ;
    LAYER M1 ;
      RECT 1595 6215 1845 9745 ;
    LAYER M1 ;
      RECT 1595 12095 1845 15625 ;
    LAYER M1 ;
      RECT 2025 335 2275 3865 ;
    LAYER M1 ;
      RECT 2025 4115 2275 5125 ;
    LAYER M1 ;
      RECT 2025 6215 2275 9745 ;
    LAYER M1 ;
      RECT 2025 9995 2275 11005 ;
    LAYER M1 ;
      RECT 2025 12095 2275 15625 ;
    LAYER M1 ;
      RECT 2025 15875 2275 16885 ;
    LAYER M1 ;
      RECT 2025 17975 2275 18985 ;
    LAYER M1 ;
      RECT 2455 335 2705 3865 ;
    LAYER M1 ;
      RECT 2455 6215 2705 9745 ;
    LAYER M1 ;
      RECT 2455 12095 2705 15625 ;
    LAYER M2 ;
      RECT 1120 280 2320 560 ;
    LAYER M2 ;
      RECT 1120 4480 2320 4760 ;
    LAYER M2 ;
      RECT 690 700 2750 980 ;
    LAYER M2 ;
      RECT 1120 6160 2320 6440 ;
    LAYER M2 ;
      RECT 1120 10360 2320 10640 ;
    LAYER M2 ;
      RECT 690 6580 2750 6860 ;
    LAYER M2 ;
      RECT 1120 12040 2320 12320 ;
    LAYER M2 ;
      RECT 1120 16240 2320 16520 ;
    LAYER M2 ;
      RECT 690 12460 2750 12740 ;
    LAYER M2 ;
      RECT 1120 18340 2320 18620 ;
    LAYER V1 ;
      RECT 1205 335 1375 505 ;
    LAYER V1 ;
      RECT 1205 4535 1375 4705 ;
    LAYER V1 ;
      RECT 1205 6215 1375 6385 ;
    LAYER V1 ;
      RECT 1205 10415 1375 10585 ;
    LAYER V1 ;
      RECT 1205 12095 1375 12265 ;
    LAYER V1 ;
      RECT 1205 16295 1375 16465 ;
    LAYER V1 ;
      RECT 1205 18395 1375 18565 ;
    LAYER V1 ;
      RECT 2065 335 2235 505 ;
    LAYER V1 ;
      RECT 2065 4535 2235 4705 ;
    LAYER V1 ;
      RECT 2065 6215 2235 6385 ;
    LAYER V1 ;
      RECT 2065 10415 2235 10585 ;
    LAYER V1 ;
      RECT 2065 12095 2235 12265 ;
    LAYER V1 ;
      RECT 2065 16295 2235 16465 ;
    LAYER V1 ;
      RECT 2065 18395 2235 18565 ;
    LAYER V1 ;
      RECT 775 755 945 925 ;
    LAYER V1 ;
      RECT 775 6635 945 6805 ;
    LAYER V1 ;
      RECT 775 12515 945 12685 ;
    LAYER V1 ;
      RECT 1635 755 1805 925 ;
    LAYER V1 ;
      RECT 1635 6635 1805 6805 ;
    LAYER V1 ;
      RECT 1635 12515 1805 12685 ;
    LAYER V1 ;
      RECT 2495 755 2665 925 ;
    LAYER V1 ;
      RECT 2495 6635 2665 6805 ;
    LAYER V1 ;
      RECT 2495 12515 2665 12685 ;
    LAYER V2 ;
      RECT 1215 345 1365 495 ;
    LAYER V2 ;
      RECT 1215 6225 1365 6375 ;
    LAYER V2 ;
      RECT 1215 12105 1365 12255 ;
    LAYER V2 ;
      RECT 1645 4545 1795 4695 ;
    LAYER V2 ;
      RECT 1645 10425 1795 10575 ;
    LAYER V2 ;
      RECT 1645 16305 1795 16455 ;
    LAYER V2 ;
      RECT 2075 765 2225 915 ;
    LAYER V2 ;
      RECT 2075 6645 2225 6795 ;
    LAYER V2 ;
      RECT 2075 12525 2225 12675 ;
    LAYER V2 ;
      RECT 2075 18405 2225 18555 ;
  END
END PMOS_S_81354572_X2_Y3
