MACRO STAGE2_INV_2661262
  ORIGIN 0 0 ;
  FOREIGN STAGE2_INV_2661262 0 0 ;
  SIZE 11.18 BY 15.12 ;
  PIN VI
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8 12.04 10.06 12.32 ;
      LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
      LAYER M2 ;
        RECT 9.3 12.04 9.62 12.32 ;
      LAYER M3 ;
        RECT 9.32 2.94 9.6 12.18 ;
      LAYER M2 ;
        RECT 9.3 2.8 9.62 3.08 ;
    END
  END VI
  PIN SN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.73 0.68 4.01 6.88 ;
      LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
      LAYER M3 ;
        RECT 3.73 6.115 4.01 6.485 ;
      LAYER M2 ;
        RECT 3.87 6.16 8.6 6.44 ;
      LAYER M3 ;
        RECT 8.46 6.115 8.74 6.485 ;
    END
  END SN
  PIN VO
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 7.84 5.76 8.12 ;
      LAYER M2 ;
        RECT 2.41 7 3.61 7.28 ;
      LAYER M2 ;
        RECT 2.85 7.84 3.17 8.12 ;
      LAYER M3 ;
        RECT 2.87 7.14 3.15 7.98 ;
      LAYER M2 ;
        RECT 2.85 7 3.17 7.28 ;
    END
  END VO
  PIN SP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.73 8.24 4.01 14.44 ;
      LAYER M3 ;
        RECT 8.46 8.24 8.74 14.44 ;
      LAYER M3 ;
        RECT 3.73 13.675 4.01 14.045 ;
      LAYER M2 ;
        RECT 3.87 13.72 8.6 14 ;
      LAYER M3 ;
        RECT 8.46 13.675 8.74 14.045 ;
    END
  END SP
  OBS 
  LAYER M2 ;
        RECT 1.12 12.04 5.76 12.32 ;
  LAYER M2 ;
        RECT 2.41 2.8 3.61 3.08 ;
  LAYER M2 ;
        RECT 8 7.84 10.06 8.12 ;
  LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 2.94 2.72 12.18 ;
  LAYER M2 ;
        RECT 2.42 2.8 2.74 3.08 ;
  LAYER M3 ;
        RECT 2.44 7.375 2.72 7.745 ;
  LAYER M2 ;
        RECT 2.58 7.42 7.31 7.7 ;
  LAYER M1 ;
        RECT 7.185 7.56 7.435 7.98 ;
  LAYER M2 ;
        RECT 7.31 7.84 8.17 8.12 ;
  LAYER M2 ;
        RECT 8.87 7.84 9.19 8.12 ;
  LAYER M3 ;
        RECT 8.89 7.14 9.17 7.98 ;
  LAYER M2 ;
        RECT 8.87 7 9.19 7.28 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 12.02 2.72 12.34 ;
  LAYER M2 ;
        RECT 2.42 2.8 2.74 3.08 ;
  LAYER M3 ;
        RECT 2.44 2.78 2.72 3.1 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 12.02 2.72 12.34 ;
  LAYER M2 ;
        RECT 2.42 2.8 2.74 3.08 ;
  LAYER M3 ;
        RECT 2.44 2.78 2.72 3.1 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.065 ;
  LAYER M2 ;
        RECT 7.14 7.84 7.48 8.12 ;
  LAYER M1 ;
        RECT 7.185 7.475 7.435 7.645 ;
  LAYER M2 ;
        RECT 7.14 7.42 7.48 7.7 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 12.02 2.72 12.34 ;
  LAYER M2 ;
        RECT 2.42 7.42 2.74 7.7 ;
  LAYER M3 ;
        RECT 2.44 7.4 2.72 7.72 ;
  LAYER M2 ;
        RECT 2.42 2.8 2.74 3.08 ;
  LAYER M3 ;
        RECT 2.44 2.78 2.72 3.1 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.065 ;
  LAYER M2 ;
        RECT 7.14 7.84 7.48 8.12 ;
  LAYER M1 ;
        RECT 7.185 7.475 7.435 7.645 ;
  LAYER M2 ;
        RECT 7.14 7.42 7.48 7.7 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 12.02 2.72 12.34 ;
  LAYER M2 ;
        RECT 2.42 7.42 2.74 7.7 ;
  LAYER M3 ;
        RECT 2.44 7.4 2.72 7.72 ;
  LAYER M2 ;
        RECT 2.42 2.8 2.74 3.08 ;
  LAYER M3 ;
        RECT 2.44 2.78 2.72 3.1 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.065 ;
  LAYER M2 ;
        RECT 7.14 7.84 7.48 8.12 ;
  LAYER M1 ;
        RECT 7.185 7.475 7.435 7.645 ;
  LAYER M2 ;
        RECT 7.14 7.42 7.48 7.7 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 12.02 2.72 12.34 ;
  LAYER M2 ;
        RECT 2.42 7.42 2.74 7.7 ;
  LAYER M3 ;
        RECT 2.44 7.4 2.72 7.72 ;
  LAYER M2 ;
        RECT 2.42 2.8 2.74 3.08 ;
  LAYER M3 ;
        RECT 2.44 2.78 2.72 3.1 ;
  LAYER M2 ;
        RECT 8.87 7.84 9.19 8.12 ;
  LAYER M3 ;
        RECT 8.89 7.82 9.17 8.14 ;
  LAYER M2 ;
        RECT 8.87 7 9.19 7.28 ;
  LAYER M3 ;
        RECT 8.89 6.98 9.17 7.3 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.065 ;
  LAYER M2 ;
        RECT 7.14 7.84 7.48 8.12 ;
  LAYER M1 ;
        RECT 7.185 7.475 7.435 7.645 ;
  LAYER M2 ;
        RECT 7.14 7.42 7.48 7.7 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 12.02 2.72 12.34 ;
  LAYER M2 ;
        RECT 2.42 7.42 2.74 7.7 ;
  LAYER M3 ;
        RECT 2.44 7.4 2.72 7.72 ;
  LAYER M2 ;
        RECT 2.42 2.8 2.74 3.08 ;
  LAYER M3 ;
        RECT 2.44 2.78 2.72 3.1 ;
  LAYER M2 ;
        RECT 8.87 7.84 9.19 8.12 ;
  LAYER M3 ;
        RECT 8.89 7.82 9.17 8.14 ;
  LAYER M2 ;
        RECT 8.87 7 9.19 7.28 ;
  LAYER M3 ;
        RECT 8.89 6.98 9.17 7.3 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M2 ;
        RECT 8.43 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 3.315 2.435 3.565 3.445 ;
  LAYER M1 ;
        RECT 3.315 0.335 3.565 1.345 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M2 ;
        RECT 2.84 6.58 4.04 6.86 ;
  LAYER M2 ;
        RECT 2.84 0.7 4.04 0.98 ;
  LAYER M2 ;
        RECT 2.41 7 3.61 7.28 ;
  LAYER M2 ;
        RECT 2.41 2.8 3.61 3.08 ;
  LAYER M3 ;
        RECT 3.73 0.68 4.01 6.88 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 14.785 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M2 ;
        RECT 7.57 8.26 10.49 8.54 ;
  LAYER M2 ;
        RECT 8 14.14 10.06 14.42 ;
  LAYER M2 ;
        RECT 8 7.84 10.06 8.12 ;
  LAYER M2 ;
        RECT 8 12.04 10.06 12.32 ;
  LAYER M3 ;
        RECT 8.46 8.24 8.74 14.44 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 11.425 ;
  LAYER M1 ;
        RECT 2.885 11.675 3.135 12.685 ;
  LAYER M1 ;
        RECT 2.885 13.775 3.135 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 11.425 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 12.685 ;
  LAYER M1 ;
        RECT 4.605 13.775 4.855 14.785 ;
  LAYER M1 ;
        RECT 5.035 7.895 5.285 11.425 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 11.425 ;
  LAYER M1 ;
        RECT 5.465 11.675 5.715 12.685 ;
  LAYER M1 ;
        RECT 5.465 13.775 5.715 14.785 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 6.19 8.54 ;
  LAYER M2 ;
        RECT 1.12 14.14 5.76 14.42 ;
  LAYER M2 ;
        RECT 1.12 7.84 5.76 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 5.76 12.32 ;
  LAYER M3 ;
        RECT 3.73 8.24 4.01 14.44 ;
  END 
END STAGE2_INV_2661262
