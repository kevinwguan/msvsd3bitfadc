* NGSPICE file created from INVERTER.ext - technology: sky130A

.subckt INVERTER vdd gate vout vss
X0 vout gate vdd vdd sky130_fd_pr__pfet_01v8 ad=2.94e+11p pd=2.66e+06u as=5.565e+11p ps=5.26e+06u w=1.05e+06u l=150000u
X1 vdd gate vout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X2 vout gate vss vss sky130_fd_pr__nfet_01v8 ad=2.94e+11p pd=2.66e+06u as=5.565e+11p ps=5.26e+06u w=1.05e+06u l=150000u
X3 vss gate vout vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
.ends

