magic
tech sky130A
magscale 1 2
timestamp 1678495828
<< nwell >>
rect 1548 1512 3268 3024
rect 860 0 3268 1512
<< pwell >>
rect 215 2718 301 2994
rect 731 2718 817 2994
rect 1247 2718 1333 2994
rect 121 1948 395 2210
rect 637 1948 911 2210
rect 1153 1948 1427 2210
rect 293 814 739 1076
rect 387 30 645 306
<< nmos >>
rect 200 1974 230 2184
rect 286 1974 316 2184
rect 716 1974 746 2184
rect 802 1974 832 2184
rect 1232 1974 1262 2184
rect 1318 1974 1348 2184
rect 372 840 402 1050
rect 458 840 488 1050
rect 544 840 574 1050
rect 630 840 660 1050
<< pmos >>
rect 1748 1974 1778 2184
rect 1834 1974 1864 2184
rect 1920 1974 1950 2184
rect 2006 1974 2036 2184
rect 2092 1974 2122 2184
rect 2178 1974 2208 2184
rect 2608 1974 2638 2184
rect 2694 1974 2724 2184
rect 2780 1974 2810 2184
rect 2866 1974 2896 2184
rect 2952 1974 2982 2184
rect 3038 1974 3068 2184
rect 1060 840 1090 1050
rect 1146 840 1176 1050
rect 1232 840 1262 1050
rect 1318 840 1348 1050
rect 1404 840 1434 1050
rect 1490 840 1520 1050
rect 1576 840 1606 1050
rect 1662 840 1692 1050
rect 1748 840 1778 1050
rect 1834 840 1864 1050
rect 1920 840 1950 1050
rect 2006 840 2036 1050
rect 2436 840 2466 1050
rect 2522 840 2552 1050
rect 2608 840 2638 1050
rect 2694 840 2724 1050
rect 2780 840 2810 1050
rect 2866 840 2896 1050
rect 2952 840 2982 1050
rect 3038 840 3068 1050
<< ndiff >>
rect 147 2160 200 2184
rect 147 2126 155 2160
rect 189 2126 200 2160
rect 147 2092 200 2126
rect 147 2058 155 2092
rect 189 2058 200 2092
rect 147 2024 200 2058
rect 147 1990 155 2024
rect 189 1990 200 2024
rect 147 1974 200 1990
rect 230 2160 286 2184
rect 230 2126 241 2160
rect 275 2126 286 2160
rect 230 2092 286 2126
rect 230 2058 241 2092
rect 275 2058 286 2092
rect 230 2024 286 2058
rect 230 1990 241 2024
rect 275 1990 286 2024
rect 230 1974 286 1990
rect 316 2160 369 2184
rect 316 2126 327 2160
rect 361 2126 369 2160
rect 316 2092 369 2126
rect 316 2058 327 2092
rect 361 2058 369 2092
rect 316 2024 369 2058
rect 316 1990 327 2024
rect 361 1990 369 2024
rect 316 1974 369 1990
rect 663 2160 716 2184
rect 663 2126 671 2160
rect 705 2126 716 2160
rect 663 2092 716 2126
rect 663 2058 671 2092
rect 705 2058 716 2092
rect 663 2024 716 2058
rect 663 1990 671 2024
rect 705 1990 716 2024
rect 663 1974 716 1990
rect 746 2160 802 2184
rect 746 2126 757 2160
rect 791 2126 802 2160
rect 746 2092 802 2126
rect 746 2058 757 2092
rect 791 2058 802 2092
rect 746 2024 802 2058
rect 746 1990 757 2024
rect 791 1990 802 2024
rect 746 1974 802 1990
rect 832 2160 885 2184
rect 832 2126 843 2160
rect 877 2126 885 2160
rect 832 2092 885 2126
rect 832 2058 843 2092
rect 877 2058 885 2092
rect 832 2024 885 2058
rect 832 1990 843 2024
rect 877 1990 885 2024
rect 832 1974 885 1990
rect 1179 2160 1232 2184
rect 1179 2126 1187 2160
rect 1221 2126 1232 2160
rect 1179 2092 1232 2126
rect 1179 2058 1187 2092
rect 1221 2058 1232 2092
rect 1179 2024 1232 2058
rect 1179 1990 1187 2024
rect 1221 1990 1232 2024
rect 1179 1974 1232 1990
rect 1262 2160 1318 2184
rect 1262 2126 1273 2160
rect 1307 2126 1318 2160
rect 1262 2092 1318 2126
rect 1262 2058 1273 2092
rect 1307 2058 1318 2092
rect 1262 2024 1318 2058
rect 1262 1990 1273 2024
rect 1307 1990 1318 2024
rect 1262 1974 1318 1990
rect 1348 2160 1401 2184
rect 1348 2126 1359 2160
rect 1393 2126 1401 2160
rect 1348 2092 1401 2126
rect 1348 2058 1359 2092
rect 1393 2058 1401 2092
rect 1348 2024 1401 2058
rect 1348 1990 1359 2024
rect 1393 1990 1401 2024
rect 1348 1974 1401 1990
rect 319 1034 372 1050
rect 319 1000 327 1034
rect 361 1000 372 1034
rect 319 966 372 1000
rect 319 932 327 966
rect 361 932 372 966
rect 319 898 372 932
rect 319 864 327 898
rect 361 864 372 898
rect 319 840 372 864
rect 402 1034 458 1050
rect 402 1000 413 1034
rect 447 1000 458 1034
rect 402 966 458 1000
rect 402 932 413 966
rect 447 932 458 966
rect 402 898 458 932
rect 402 864 413 898
rect 447 864 458 898
rect 402 840 458 864
rect 488 1034 544 1050
rect 488 1000 499 1034
rect 533 1000 544 1034
rect 488 966 544 1000
rect 488 932 499 966
rect 533 932 544 966
rect 488 898 544 932
rect 488 864 499 898
rect 533 864 544 898
rect 488 840 544 864
rect 574 1034 630 1050
rect 574 1000 585 1034
rect 619 1000 630 1034
rect 574 966 630 1000
rect 574 932 585 966
rect 619 932 630 966
rect 574 898 630 932
rect 574 864 585 898
rect 619 864 630 898
rect 574 840 630 864
rect 660 1034 713 1050
rect 660 1000 671 1034
rect 705 1000 713 1034
rect 660 966 713 1000
rect 660 932 671 966
rect 705 932 713 966
rect 660 898 713 932
rect 660 864 671 898
rect 705 864 713 898
rect 660 840 713 864
<< pdiff >>
rect 1695 2160 1748 2184
rect 1695 2126 1703 2160
rect 1737 2126 1748 2160
rect 1695 2092 1748 2126
rect 1695 2058 1703 2092
rect 1737 2058 1748 2092
rect 1695 2024 1748 2058
rect 1695 1990 1703 2024
rect 1737 1990 1748 2024
rect 1695 1974 1748 1990
rect 1778 2160 1834 2184
rect 1778 2126 1789 2160
rect 1823 2126 1834 2160
rect 1778 2092 1834 2126
rect 1778 2058 1789 2092
rect 1823 2058 1834 2092
rect 1778 2024 1834 2058
rect 1778 1990 1789 2024
rect 1823 1990 1834 2024
rect 1778 1974 1834 1990
rect 1864 2160 1920 2184
rect 1864 2126 1875 2160
rect 1909 2126 1920 2160
rect 1864 2092 1920 2126
rect 1864 2058 1875 2092
rect 1909 2058 1920 2092
rect 1864 2024 1920 2058
rect 1864 1990 1875 2024
rect 1909 1990 1920 2024
rect 1864 1974 1920 1990
rect 1950 2160 2006 2184
rect 1950 2126 1961 2160
rect 1995 2126 2006 2160
rect 1950 2092 2006 2126
rect 1950 2058 1961 2092
rect 1995 2058 2006 2092
rect 1950 2024 2006 2058
rect 1950 1990 1961 2024
rect 1995 1990 2006 2024
rect 1950 1974 2006 1990
rect 2036 2160 2092 2184
rect 2036 2126 2047 2160
rect 2081 2126 2092 2160
rect 2036 2092 2092 2126
rect 2036 2058 2047 2092
rect 2081 2058 2092 2092
rect 2036 2024 2092 2058
rect 2036 1990 2047 2024
rect 2081 1990 2092 2024
rect 2036 1974 2092 1990
rect 2122 2160 2178 2184
rect 2122 2126 2133 2160
rect 2167 2126 2178 2160
rect 2122 2092 2178 2126
rect 2122 2058 2133 2092
rect 2167 2058 2178 2092
rect 2122 2024 2178 2058
rect 2122 1990 2133 2024
rect 2167 1990 2178 2024
rect 2122 1974 2178 1990
rect 2208 2160 2261 2184
rect 2208 2126 2219 2160
rect 2253 2126 2261 2160
rect 2208 2092 2261 2126
rect 2208 2058 2219 2092
rect 2253 2058 2261 2092
rect 2208 2024 2261 2058
rect 2208 1990 2219 2024
rect 2253 1990 2261 2024
rect 2208 1974 2261 1990
rect 2555 2160 2608 2184
rect 2555 2126 2563 2160
rect 2597 2126 2608 2160
rect 2555 2092 2608 2126
rect 2555 2058 2563 2092
rect 2597 2058 2608 2092
rect 2555 2024 2608 2058
rect 2555 1990 2563 2024
rect 2597 1990 2608 2024
rect 2555 1974 2608 1990
rect 2638 2160 2694 2184
rect 2638 2126 2649 2160
rect 2683 2126 2694 2160
rect 2638 2092 2694 2126
rect 2638 2058 2649 2092
rect 2683 2058 2694 2092
rect 2638 2024 2694 2058
rect 2638 1990 2649 2024
rect 2683 1990 2694 2024
rect 2638 1974 2694 1990
rect 2724 2160 2780 2184
rect 2724 2126 2735 2160
rect 2769 2126 2780 2160
rect 2724 2092 2780 2126
rect 2724 2058 2735 2092
rect 2769 2058 2780 2092
rect 2724 2024 2780 2058
rect 2724 1990 2735 2024
rect 2769 1990 2780 2024
rect 2724 1974 2780 1990
rect 2810 2160 2866 2184
rect 2810 2126 2821 2160
rect 2855 2126 2866 2160
rect 2810 2092 2866 2126
rect 2810 2058 2821 2092
rect 2855 2058 2866 2092
rect 2810 2024 2866 2058
rect 2810 1990 2821 2024
rect 2855 1990 2866 2024
rect 2810 1974 2866 1990
rect 2896 2160 2952 2184
rect 2896 2126 2907 2160
rect 2941 2126 2952 2160
rect 2896 2092 2952 2126
rect 2896 2058 2907 2092
rect 2941 2058 2952 2092
rect 2896 2024 2952 2058
rect 2896 1990 2907 2024
rect 2941 1990 2952 2024
rect 2896 1974 2952 1990
rect 2982 2160 3038 2184
rect 2982 2126 2993 2160
rect 3027 2126 3038 2160
rect 2982 2092 3038 2126
rect 2982 2058 2993 2092
rect 3027 2058 3038 2092
rect 2982 2024 3038 2058
rect 2982 1990 2993 2024
rect 3027 1990 3038 2024
rect 2982 1974 3038 1990
rect 3068 2160 3121 2184
rect 3068 2126 3079 2160
rect 3113 2126 3121 2160
rect 3068 2092 3121 2126
rect 3068 2058 3079 2092
rect 3113 2058 3121 2092
rect 3068 2024 3121 2058
rect 3068 1990 3079 2024
rect 3113 1990 3121 2024
rect 3068 1974 3121 1990
rect 1007 1034 1060 1050
rect 1007 1000 1015 1034
rect 1049 1000 1060 1034
rect 1007 966 1060 1000
rect 1007 932 1015 966
rect 1049 932 1060 966
rect 1007 898 1060 932
rect 1007 864 1015 898
rect 1049 864 1060 898
rect 1007 840 1060 864
rect 1090 1034 1146 1050
rect 1090 1000 1101 1034
rect 1135 1000 1146 1034
rect 1090 966 1146 1000
rect 1090 932 1101 966
rect 1135 932 1146 966
rect 1090 898 1146 932
rect 1090 864 1101 898
rect 1135 864 1146 898
rect 1090 840 1146 864
rect 1176 1034 1232 1050
rect 1176 1000 1187 1034
rect 1221 1000 1232 1034
rect 1176 966 1232 1000
rect 1176 932 1187 966
rect 1221 932 1232 966
rect 1176 898 1232 932
rect 1176 864 1187 898
rect 1221 864 1232 898
rect 1176 840 1232 864
rect 1262 1034 1318 1050
rect 1262 1000 1273 1034
rect 1307 1000 1318 1034
rect 1262 966 1318 1000
rect 1262 932 1273 966
rect 1307 932 1318 966
rect 1262 898 1318 932
rect 1262 864 1273 898
rect 1307 864 1318 898
rect 1262 840 1318 864
rect 1348 1034 1404 1050
rect 1348 1000 1359 1034
rect 1393 1000 1404 1034
rect 1348 966 1404 1000
rect 1348 932 1359 966
rect 1393 932 1404 966
rect 1348 898 1404 932
rect 1348 864 1359 898
rect 1393 864 1404 898
rect 1348 840 1404 864
rect 1434 1034 1490 1050
rect 1434 1000 1445 1034
rect 1479 1000 1490 1034
rect 1434 966 1490 1000
rect 1434 932 1445 966
rect 1479 932 1490 966
rect 1434 898 1490 932
rect 1434 864 1445 898
rect 1479 864 1490 898
rect 1434 840 1490 864
rect 1520 1034 1576 1050
rect 1520 1000 1531 1034
rect 1565 1000 1576 1034
rect 1520 966 1576 1000
rect 1520 932 1531 966
rect 1565 932 1576 966
rect 1520 898 1576 932
rect 1520 864 1531 898
rect 1565 864 1576 898
rect 1520 840 1576 864
rect 1606 1034 1662 1050
rect 1606 1000 1617 1034
rect 1651 1000 1662 1034
rect 1606 966 1662 1000
rect 1606 932 1617 966
rect 1651 932 1662 966
rect 1606 898 1662 932
rect 1606 864 1617 898
rect 1651 864 1662 898
rect 1606 840 1662 864
rect 1692 1034 1748 1050
rect 1692 1000 1703 1034
rect 1737 1000 1748 1034
rect 1692 966 1748 1000
rect 1692 932 1703 966
rect 1737 932 1748 966
rect 1692 898 1748 932
rect 1692 864 1703 898
rect 1737 864 1748 898
rect 1692 840 1748 864
rect 1778 1034 1834 1050
rect 1778 1000 1789 1034
rect 1823 1000 1834 1034
rect 1778 966 1834 1000
rect 1778 932 1789 966
rect 1823 932 1834 966
rect 1778 898 1834 932
rect 1778 864 1789 898
rect 1823 864 1834 898
rect 1778 840 1834 864
rect 1864 1034 1920 1050
rect 1864 1000 1875 1034
rect 1909 1000 1920 1034
rect 1864 966 1920 1000
rect 1864 932 1875 966
rect 1909 932 1920 966
rect 1864 898 1920 932
rect 1864 864 1875 898
rect 1909 864 1920 898
rect 1864 840 1920 864
rect 1950 1034 2006 1050
rect 1950 1000 1961 1034
rect 1995 1000 2006 1034
rect 1950 966 2006 1000
rect 1950 932 1961 966
rect 1995 932 2006 966
rect 1950 898 2006 932
rect 1950 864 1961 898
rect 1995 864 2006 898
rect 1950 840 2006 864
rect 2036 1034 2089 1050
rect 2036 1000 2047 1034
rect 2081 1000 2089 1034
rect 2036 966 2089 1000
rect 2036 932 2047 966
rect 2081 932 2089 966
rect 2036 898 2089 932
rect 2036 864 2047 898
rect 2081 864 2089 898
rect 2036 840 2089 864
rect 2383 1034 2436 1050
rect 2383 1000 2391 1034
rect 2425 1000 2436 1034
rect 2383 966 2436 1000
rect 2383 932 2391 966
rect 2425 932 2436 966
rect 2383 898 2436 932
rect 2383 864 2391 898
rect 2425 864 2436 898
rect 2383 840 2436 864
rect 2466 1034 2522 1050
rect 2466 1000 2477 1034
rect 2511 1000 2522 1034
rect 2466 966 2522 1000
rect 2466 932 2477 966
rect 2511 932 2522 966
rect 2466 898 2522 932
rect 2466 864 2477 898
rect 2511 864 2522 898
rect 2466 840 2522 864
rect 2552 1034 2608 1050
rect 2552 1000 2563 1034
rect 2597 1000 2608 1034
rect 2552 966 2608 1000
rect 2552 932 2563 966
rect 2597 932 2608 966
rect 2552 898 2608 932
rect 2552 864 2563 898
rect 2597 864 2608 898
rect 2552 840 2608 864
rect 2638 1034 2694 1050
rect 2638 1000 2649 1034
rect 2683 1000 2694 1034
rect 2638 966 2694 1000
rect 2638 932 2649 966
rect 2683 932 2694 966
rect 2638 898 2694 932
rect 2638 864 2649 898
rect 2683 864 2694 898
rect 2638 840 2694 864
rect 2724 1034 2780 1050
rect 2724 1000 2735 1034
rect 2769 1000 2780 1034
rect 2724 966 2780 1000
rect 2724 932 2735 966
rect 2769 932 2780 966
rect 2724 898 2780 932
rect 2724 864 2735 898
rect 2769 864 2780 898
rect 2724 840 2780 864
rect 2810 1034 2866 1050
rect 2810 1000 2821 1034
rect 2855 1000 2866 1034
rect 2810 966 2866 1000
rect 2810 932 2821 966
rect 2855 932 2866 966
rect 2810 898 2866 932
rect 2810 864 2821 898
rect 2855 864 2866 898
rect 2810 840 2866 864
rect 2896 1034 2952 1050
rect 2896 1000 2907 1034
rect 2941 1000 2952 1034
rect 2896 966 2952 1000
rect 2896 932 2907 966
rect 2941 932 2952 966
rect 2896 898 2952 932
rect 2896 864 2907 898
rect 2941 864 2952 898
rect 2896 840 2952 864
rect 2982 1034 3038 1050
rect 2982 1000 2993 1034
rect 3027 1000 3038 1034
rect 2982 966 3038 1000
rect 2982 932 2993 966
rect 3027 932 3038 966
rect 2982 898 3038 932
rect 2982 864 2993 898
rect 3027 864 3038 898
rect 2982 840 3038 864
rect 3068 1034 3121 1050
rect 3068 1000 3079 1034
rect 3113 1000 3121 1034
rect 3068 966 3121 1000
rect 3068 932 3079 966
rect 3113 932 3121 966
rect 3068 898 3121 932
rect 3068 864 3079 898
rect 3113 864 3121 898
rect 3068 840 3121 864
<< ndiffc >>
rect 155 2126 189 2160
rect 155 2058 189 2092
rect 155 1990 189 2024
rect 241 2126 275 2160
rect 241 2058 275 2092
rect 241 1990 275 2024
rect 327 2126 361 2160
rect 327 2058 361 2092
rect 327 1990 361 2024
rect 671 2126 705 2160
rect 671 2058 705 2092
rect 671 1990 705 2024
rect 757 2126 791 2160
rect 757 2058 791 2092
rect 757 1990 791 2024
rect 843 2126 877 2160
rect 843 2058 877 2092
rect 843 1990 877 2024
rect 1187 2126 1221 2160
rect 1187 2058 1221 2092
rect 1187 1990 1221 2024
rect 1273 2126 1307 2160
rect 1273 2058 1307 2092
rect 1273 1990 1307 2024
rect 1359 2126 1393 2160
rect 1359 2058 1393 2092
rect 1359 1990 1393 2024
rect 327 1000 361 1034
rect 327 932 361 966
rect 327 864 361 898
rect 413 1000 447 1034
rect 413 932 447 966
rect 413 864 447 898
rect 499 1000 533 1034
rect 499 932 533 966
rect 499 864 533 898
rect 585 1000 619 1034
rect 585 932 619 966
rect 585 864 619 898
rect 671 1000 705 1034
rect 671 932 705 966
rect 671 864 705 898
<< pdiffc >>
rect 1703 2126 1737 2160
rect 1703 2058 1737 2092
rect 1703 1990 1737 2024
rect 1789 2126 1823 2160
rect 1789 2058 1823 2092
rect 1789 1990 1823 2024
rect 1875 2126 1909 2160
rect 1875 2058 1909 2092
rect 1875 1990 1909 2024
rect 1961 2126 1995 2160
rect 1961 2058 1995 2092
rect 1961 1990 1995 2024
rect 2047 2126 2081 2160
rect 2047 2058 2081 2092
rect 2047 1990 2081 2024
rect 2133 2126 2167 2160
rect 2133 2058 2167 2092
rect 2133 1990 2167 2024
rect 2219 2126 2253 2160
rect 2219 2058 2253 2092
rect 2219 1990 2253 2024
rect 2563 2126 2597 2160
rect 2563 2058 2597 2092
rect 2563 1990 2597 2024
rect 2649 2126 2683 2160
rect 2649 2058 2683 2092
rect 2649 1990 2683 2024
rect 2735 2126 2769 2160
rect 2735 2058 2769 2092
rect 2735 1990 2769 2024
rect 2821 2126 2855 2160
rect 2821 2058 2855 2092
rect 2821 1990 2855 2024
rect 2907 2126 2941 2160
rect 2907 2058 2941 2092
rect 2907 1990 2941 2024
rect 2993 2126 3027 2160
rect 2993 2058 3027 2092
rect 2993 1990 3027 2024
rect 3079 2126 3113 2160
rect 3079 2058 3113 2092
rect 3079 1990 3113 2024
rect 1015 1000 1049 1034
rect 1015 932 1049 966
rect 1015 864 1049 898
rect 1101 1000 1135 1034
rect 1101 932 1135 966
rect 1101 864 1135 898
rect 1187 1000 1221 1034
rect 1187 932 1221 966
rect 1187 864 1221 898
rect 1273 1000 1307 1034
rect 1273 932 1307 966
rect 1273 864 1307 898
rect 1359 1000 1393 1034
rect 1359 932 1393 966
rect 1359 864 1393 898
rect 1445 1000 1479 1034
rect 1445 932 1479 966
rect 1445 864 1479 898
rect 1531 1000 1565 1034
rect 1531 932 1565 966
rect 1531 864 1565 898
rect 1617 1000 1651 1034
rect 1617 932 1651 966
rect 1617 864 1651 898
rect 1703 1000 1737 1034
rect 1703 932 1737 966
rect 1703 864 1737 898
rect 1789 1000 1823 1034
rect 1789 932 1823 966
rect 1789 864 1823 898
rect 1875 1000 1909 1034
rect 1875 932 1909 966
rect 1875 864 1909 898
rect 1961 1000 1995 1034
rect 1961 932 1995 966
rect 1961 864 1995 898
rect 2047 1000 2081 1034
rect 2047 932 2081 966
rect 2047 864 2081 898
rect 2391 1000 2425 1034
rect 2391 932 2425 966
rect 2391 864 2425 898
rect 2477 1000 2511 1034
rect 2477 932 2511 966
rect 2477 864 2511 898
rect 2563 1000 2597 1034
rect 2563 932 2597 966
rect 2563 864 2597 898
rect 2649 1000 2683 1034
rect 2649 932 2683 966
rect 2649 864 2683 898
rect 2735 1000 2769 1034
rect 2735 932 2769 966
rect 2735 864 2769 898
rect 2821 1000 2855 1034
rect 2821 932 2855 966
rect 2821 864 2855 898
rect 2907 1000 2941 1034
rect 2907 932 2941 966
rect 2907 864 2941 898
rect 2993 1000 3027 1034
rect 2993 932 3027 966
rect 2993 864 3027 898
rect 3079 1000 3113 1034
rect 3079 932 3113 966
rect 3079 864 3113 898
<< psubdiff >>
rect 241 2873 275 2968
rect 241 2744 275 2839
rect 757 2873 791 2968
rect 757 2744 791 2839
rect 1273 2873 1307 2968
rect 1273 2744 1307 2839
rect 413 185 447 280
rect 413 56 447 151
rect 585 185 619 280
rect 585 56 619 151
<< nsubdiff >>
rect 1789 2873 1823 2968
rect 1789 2744 1823 2839
rect 1961 2873 1995 2968
rect 1961 2744 1995 2839
rect 2133 2873 2167 2968
rect 2133 2744 2167 2839
rect 2649 2873 2683 2968
rect 2649 2744 2683 2839
rect 2821 2873 2855 2968
rect 2821 2744 2855 2839
rect 2993 2873 3027 2968
rect 2993 2744 3027 2839
rect 1101 185 1135 280
rect 1101 56 1135 151
rect 1273 185 1307 280
rect 1273 56 1307 151
rect 1445 185 1479 280
rect 1445 56 1479 151
rect 1617 185 1651 280
rect 1617 56 1651 151
rect 1789 185 1823 280
rect 1789 56 1823 151
rect 1961 185 1995 280
rect 1961 56 1995 151
rect 2477 185 2511 280
rect 2477 56 2511 151
rect 2649 185 2683 280
rect 2649 56 2683 151
rect 2821 185 2855 280
rect 2821 56 2855 151
rect 2993 185 3027 280
rect 2993 56 3027 151
<< psubdiffcont >>
rect 241 2839 275 2873
rect 757 2839 791 2873
rect 1273 2839 1307 2873
rect 413 151 447 185
rect 585 151 619 185
<< nsubdiffcont >>
rect 1789 2839 1823 2873
rect 1961 2839 1995 2873
rect 2133 2839 2167 2873
rect 2649 2839 2683 2873
rect 2821 2839 2855 2873
rect 2993 2839 3027 2873
rect 1101 151 1135 185
rect 1273 151 1307 185
rect 1445 151 1479 185
rect 1617 151 1651 185
rect 1789 151 1823 185
rect 1961 151 1995 185
rect 2477 151 2511 185
rect 2649 151 2683 185
rect 2821 151 2855 185
rect 2993 151 3027 185
<< poly >>
rect 200 2453 316 2463
rect 200 2419 241 2453
rect 275 2419 316 2453
rect 200 2409 316 2419
rect 200 2184 230 2409
rect 286 2184 316 2409
rect 716 2453 832 2463
rect 716 2419 757 2453
rect 791 2419 832 2453
rect 716 2409 832 2419
rect 716 2184 746 2409
rect 802 2184 832 2409
rect 1232 2453 1348 2463
rect 1232 2419 1273 2453
rect 1307 2419 1348 2453
rect 1232 2409 1348 2419
rect 1232 2184 1262 2409
rect 1318 2184 1348 2409
rect 1748 2453 1864 2463
rect 1748 2419 1789 2453
rect 1823 2419 1864 2453
rect 1748 2409 1864 2419
rect 1748 2184 1778 2409
rect 1834 2184 1864 2409
rect 1920 2453 2036 2463
rect 1920 2419 1961 2453
rect 1995 2419 2036 2453
rect 1920 2409 2036 2419
rect 1920 2184 1950 2409
rect 2006 2184 2036 2409
rect 2092 2453 2208 2463
rect 2092 2419 2133 2453
rect 2167 2419 2208 2453
rect 2092 2409 2208 2419
rect 2092 2184 2122 2409
rect 2178 2184 2208 2409
rect 2608 2453 2724 2463
rect 2608 2419 2649 2453
rect 2683 2419 2724 2453
rect 2608 2409 2724 2419
rect 2608 2184 2638 2409
rect 2694 2184 2724 2409
rect 2780 2453 2896 2463
rect 2780 2419 2821 2453
rect 2855 2419 2896 2453
rect 2780 2409 2896 2419
rect 2780 2184 2810 2409
rect 2866 2184 2896 2409
rect 2952 2453 3068 2463
rect 2952 2419 2993 2453
rect 3027 2419 3068 2453
rect 2952 2409 3068 2419
rect 2952 2184 2982 2409
rect 3038 2184 3068 2409
rect 200 1764 230 1974
rect 286 1764 316 1974
rect 716 1764 746 1974
rect 802 1764 832 1974
rect 1232 1764 1262 1974
rect 1318 1764 1348 1974
rect 1748 1764 1778 1974
rect 1834 1764 1864 1974
rect 1920 1764 1950 1974
rect 2006 1764 2036 1974
rect 2092 1764 2122 1974
rect 2178 1764 2208 1974
rect 2608 1764 2638 1974
rect 2694 1764 2724 1974
rect 2780 1764 2810 1974
rect 2866 1764 2896 1974
rect 2952 1764 2982 1974
rect 3038 1764 3068 1974
rect 372 1050 402 1260
rect 458 1050 488 1260
rect 544 1050 574 1260
rect 630 1050 660 1260
rect 1060 1050 1090 1260
rect 1146 1050 1176 1260
rect 1232 1050 1262 1260
rect 1318 1050 1348 1260
rect 1404 1050 1434 1260
rect 1490 1050 1520 1260
rect 1576 1050 1606 1260
rect 1662 1050 1692 1260
rect 1748 1050 1778 1260
rect 1834 1050 1864 1260
rect 1920 1050 1950 1260
rect 2006 1050 2036 1260
rect 2436 1050 2466 1260
rect 2522 1050 2552 1260
rect 2608 1050 2638 1260
rect 2694 1050 2724 1260
rect 2780 1050 2810 1260
rect 2866 1050 2896 1260
rect 2952 1050 2982 1260
rect 3038 1050 3068 1260
rect 372 615 402 840
rect 458 615 488 840
rect 372 605 488 615
rect 372 571 413 605
rect 447 571 488 605
rect 372 561 488 571
rect 544 615 574 840
rect 630 615 660 840
rect 544 605 660 615
rect 544 571 585 605
rect 619 571 660 605
rect 544 561 660 571
rect 1060 615 1090 840
rect 1146 615 1176 840
rect 1060 605 1176 615
rect 1060 571 1101 605
rect 1135 571 1176 605
rect 1060 561 1176 571
rect 1232 615 1262 840
rect 1318 615 1348 840
rect 1232 605 1348 615
rect 1232 571 1273 605
rect 1307 571 1348 605
rect 1232 561 1348 571
rect 1404 615 1434 840
rect 1490 615 1520 840
rect 1404 605 1520 615
rect 1404 571 1445 605
rect 1479 571 1520 605
rect 1404 561 1520 571
rect 1576 615 1606 840
rect 1662 615 1692 840
rect 1576 605 1692 615
rect 1576 571 1617 605
rect 1651 571 1692 605
rect 1576 561 1692 571
rect 1748 615 1778 840
rect 1834 615 1864 840
rect 1748 605 1864 615
rect 1748 571 1789 605
rect 1823 571 1864 605
rect 1748 561 1864 571
rect 1920 615 1950 840
rect 2006 615 2036 840
rect 1920 605 2036 615
rect 1920 571 1961 605
rect 1995 571 2036 605
rect 1920 561 2036 571
rect 2436 615 2466 840
rect 2522 615 2552 840
rect 2436 605 2552 615
rect 2436 571 2477 605
rect 2511 571 2552 605
rect 2436 561 2552 571
rect 2608 615 2638 840
rect 2694 615 2724 840
rect 2608 605 2724 615
rect 2608 571 2649 605
rect 2683 571 2724 605
rect 2608 561 2724 571
rect 2780 615 2810 840
rect 2866 615 2896 840
rect 2780 605 2896 615
rect 2780 571 2821 605
rect 2855 571 2896 605
rect 2780 561 2896 571
rect 2952 615 2982 840
rect 3038 615 3068 840
rect 2952 605 3068 615
rect 2952 571 2993 605
rect 3027 571 3068 605
rect 2952 561 3068 571
<< polycont >>
rect 241 2419 275 2453
rect 757 2419 791 2453
rect 1273 2419 1307 2453
rect 1789 2419 1823 2453
rect 1961 2419 1995 2453
rect 2133 2419 2167 2453
rect 2649 2419 2683 2453
rect 2821 2419 2855 2453
rect 2993 2419 3027 2453
rect 413 571 447 605
rect 585 571 619 605
rect 1101 571 1135 605
rect 1273 571 1307 605
rect 1445 571 1479 605
rect 1617 571 1651 605
rect 1789 571 1823 605
rect 1961 571 1995 605
rect 2477 571 2511 605
rect 2649 571 2683 605
rect 2821 571 2855 605
rect 2993 571 3027 605
<< locali >>
rect 233 2873 283 2957
rect 749 2873 799 2957
rect 233 2839 241 2873
rect 275 2839 283 2873
rect 233 2755 283 2839
rect 405 2839 413 2873
rect 447 2839 455 2873
rect 405 2789 455 2839
rect 405 2755 413 2789
rect 447 2755 455 2789
rect 749 2839 757 2873
rect 791 2839 799 2873
rect 749 2755 799 2839
rect 1265 2873 1315 2957
rect 1265 2839 1273 2873
rect 1307 2839 1315 2873
rect 1265 2755 1315 2839
rect 1781 2873 1831 2957
rect 1781 2839 1789 2873
rect 1823 2839 1831 2873
rect 1781 2755 1831 2839
rect 1953 2873 2003 2957
rect 1953 2839 1961 2873
rect 1995 2839 2003 2873
rect 1953 2755 2003 2839
rect 2125 2873 2175 2957
rect 2125 2839 2133 2873
rect 2167 2839 2175 2873
rect 2125 2755 2175 2839
rect 2641 2873 2691 2957
rect 2641 2839 2649 2873
rect 2683 2839 2691 2873
rect 2641 2755 2691 2839
rect 2813 2873 2863 2957
rect 2813 2839 2821 2873
rect 2855 2839 2863 2873
rect 2813 2755 2863 2839
rect 2985 2873 3035 2957
rect 2985 2839 2993 2873
rect 3027 2839 3035 2873
rect 2985 2755 3035 2839
rect 233 2453 283 2537
rect 233 2419 241 2453
rect 275 2419 283 2453
rect 233 2335 283 2419
rect 749 2453 799 2537
rect 749 2419 757 2453
rect 791 2419 799 2453
rect 749 2335 799 2419
rect 1265 2453 1315 2537
rect 1781 2453 1831 2537
rect 1265 2419 1273 2453
rect 1307 2419 1315 2453
rect 1265 2335 1315 2419
rect 1695 2419 1703 2453
rect 1737 2419 1745 2453
rect 1695 2369 1745 2419
rect 1695 2335 1703 2369
rect 1737 2335 1745 2369
rect 1781 2419 1789 2453
rect 1823 2419 1831 2453
rect 1781 2335 1831 2419
rect 1953 2453 2003 2537
rect 1953 2419 1961 2453
rect 1995 2419 2003 2453
rect 1953 2335 2003 2419
rect 2125 2453 2175 2537
rect 2125 2419 2133 2453
rect 2167 2419 2175 2453
rect 2125 2335 2175 2419
rect 2641 2453 2691 2537
rect 2641 2419 2649 2453
rect 2683 2419 2691 2453
rect 2641 2335 2691 2419
rect 2813 2453 2863 2537
rect 2813 2419 2821 2453
rect 2855 2419 2863 2453
rect 2813 2335 2863 2419
rect 2985 2453 3035 2537
rect 2985 2419 2993 2453
rect 3027 2419 3035 2453
rect 2985 2335 3035 2419
rect 147 2160 197 2285
rect 147 2126 155 2160
rect 189 2126 197 2160
rect 147 2092 197 2126
rect 147 2058 155 2092
rect 189 2058 197 2092
rect 147 2024 197 2058
rect 147 1990 155 2024
rect 189 1990 197 2024
rect 147 1697 197 1990
rect 147 1663 155 1697
rect 189 1663 197 1697
rect 147 1579 197 1663
rect 233 2160 283 2285
rect 233 2126 241 2160
rect 275 2126 283 2160
rect 233 2092 283 2126
rect 233 2058 241 2092
rect 275 2058 283 2092
rect 233 2024 283 2058
rect 233 1990 241 2024
rect 275 1990 283 2024
rect 233 1613 283 1990
rect 233 1579 241 1613
rect 275 1579 283 1613
rect 319 2160 369 2285
rect 319 2126 327 2160
rect 361 2126 369 2160
rect 319 2092 369 2126
rect 319 2058 327 2092
rect 361 2058 369 2092
rect 319 2024 369 2058
rect 319 1990 327 2024
rect 361 1990 369 2024
rect 319 1697 369 1990
rect 319 1663 327 1697
rect 361 1663 369 1697
rect 319 1579 369 1663
rect 663 2160 713 2285
rect 663 2126 671 2160
rect 705 2126 713 2160
rect 663 2092 713 2126
rect 663 2058 671 2092
rect 705 2058 713 2092
rect 663 2024 713 2058
rect 663 1990 671 2024
rect 705 1990 713 2024
rect 663 1697 713 1990
rect 663 1663 671 1697
rect 705 1663 713 1697
rect 577 1579 585 1613
rect 619 1579 627 1613
rect 663 1579 713 1663
rect 749 2160 799 2285
rect 749 2126 757 2160
rect 791 2126 799 2160
rect 749 2092 799 2126
rect 749 2058 757 2092
rect 791 2058 799 2092
rect 749 2024 799 2058
rect 749 1990 757 2024
rect 791 1990 799 2024
rect 749 1613 799 1990
rect 749 1579 757 1613
rect 791 1579 799 1613
rect 835 2160 885 2285
rect 835 2126 843 2160
rect 877 2126 885 2160
rect 835 2092 885 2126
rect 835 2058 843 2092
rect 877 2058 885 2092
rect 835 2024 885 2058
rect 835 1990 843 2024
rect 877 1990 885 2024
rect 835 1697 885 1990
rect 835 1663 843 1697
rect 877 1663 885 1697
rect 835 1579 885 1663
rect 1179 2160 1229 2285
rect 1179 2126 1187 2160
rect 1221 2126 1229 2160
rect 1179 2092 1229 2126
rect 1179 2058 1187 2092
rect 1221 2058 1229 2092
rect 1179 2024 1229 2058
rect 1179 1990 1187 2024
rect 1221 1990 1229 2024
rect 1179 1697 1229 1990
rect 1179 1663 1187 1697
rect 1221 1663 1229 1697
rect 921 1579 929 1613
rect 963 1579 971 1613
rect 1179 1579 1229 1663
rect 1265 2160 1315 2285
rect 1265 2126 1273 2160
rect 1307 2126 1315 2160
rect 1265 2092 1315 2126
rect 1265 2058 1273 2092
rect 1307 2058 1315 2092
rect 1265 2024 1315 2058
rect 1265 1990 1273 2024
rect 1307 1990 1315 2024
rect 1265 1613 1315 1990
rect 1265 1579 1273 1613
rect 1307 1579 1315 1613
rect 1351 2160 1401 2285
rect 1351 2126 1359 2160
rect 1393 2126 1401 2160
rect 1351 2092 1401 2126
rect 1351 2058 1359 2092
rect 1393 2058 1401 2092
rect 1351 2024 1401 2058
rect 1351 1990 1359 2024
rect 1393 1990 1401 2024
rect 1351 1697 1401 1990
rect 1351 1663 1359 1697
rect 1393 1663 1401 1697
rect 1351 1579 1401 1663
rect 1695 2160 1745 2285
rect 1695 2126 1703 2160
rect 1737 2126 1745 2160
rect 1695 2092 1745 2126
rect 1695 2058 1703 2092
rect 1737 2058 1745 2092
rect 1695 2024 1745 2058
rect 1695 1990 1703 2024
rect 1737 1990 1745 2024
rect 1695 1697 1745 1990
rect 1695 1663 1703 1697
rect 1737 1663 1745 1697
rect 1695 1579 1745 1663
rect 1781 2160 1831 2285
rect 1781 2126 1789 2160
rect 1823 2126 1831 2160
rect 1781 2092 1831 2126
rect 1781 2058 1789 2092
rect 1823 2058 1831 2092
rect 1781 2024 1831 2058
rect 1781 1990 1789 2024
rect 1823 1990 1831 2024
rect 1781 1613 1831 1990
rect 1781 1579 1789 1613
rect 1823 1579 1831 1613
rect 1867 2160 1917 2285
rect 1867 2126 1875 2160
rect 1909 2126 1917 2160
rect 1867 2092 1917 2126
rect 1867 2058 1875 2092
rect 1909 2058 1917 2092
rect 1867 2024 1917 2058
rect 1867 1990 1875 2024
rect 1909 1990 1917 2024
rect 1867 1697 1917 1990
rect 1867 1663 1875 1697
rect 1909 1663 1917 1697
rect 1867 1579 1917 1663
rect 1953 2160 2003 2285
rect 1953 2126 1961 2160
rect 1995 2126 2003 2160
rect 1953 2092 2003 2126
rect 1953 2058 1961 2092
rect 1995 2058 2003 2092
rect 1953 2024 2003 2058
rect 1953 1990 1961 2024
rect 1995 1990 2003 2024
rect 1953 1613 2003 1990
rect 1953 1579 1961 1613
rect 1995 1579 2003 1613
rect 2039 2160 2089 2285
rect 2039 2126 2047 2160
rect 2081 2126 2089 2160
rect 2039 2092 2089 2126
rect 2039 2058 2047 2092
rect 2081 2058 2089 2092
rect 2039 2024 2089 2058
rect 2039 1990 2047 2024
rect 2081 1990 2089 2024
rect 2039 1697 2089 1990
rect 2039 1663 2047 1697
rect 2081 1663 2089 1697
rect 2039 1579 2089 1663
rect 2125 2160 2175 2285
rect 2125 2126 2133 2160
rect 2167 2126 2175 2160
rect 2125 2092 2175 2126
rect 2125 2058 2133 2092
rect 2167 2058 2175 2092
rect 2125 2024 2175 2058
rect 2125 1990 2133 2024
rect 2167 1990 2175 2024
rect 2125 1613 2175 1990
rect 2125 1579 2133 1613
rect 2167 1579 2175 1613
rect 2211 2160 2261 2285
rect 2211 2126 2219 2160
rect 2253 2126 2261 2160
rect 2211 2092 2261 2126
rect 2211 2058 2219 2092
rect 2253 2058 2261 2092
rect 2211 2024 2261 2058
rect 2211 1990 2219 2024
rect 2253 1990 2261 2024
rect 2211 1697 2261 1990
rect 2211 1663 2219 1697
rect 2253 1663 2261 1697
rect 2211 1579 2261 1663
rect 2555 2160 2605 2285
rect 2555 2126 2563 2160
rect 2597 2126 2605 2160
rect 2555 2092 2605 2126
rect 2555 2058 2563 2092
rect 2597 2058 2605 2092
rect 2555 2024 2605 2058
rect 2555 1990 2563 2024
rect 2597 1990 2605 2024
rect 2555 1697 2605 1990
rect 2555 1663 2563 1697
rect 2597 1663 2605 1697
rect 2469 1579 2477 1613
rect 2511 1579 2519 1613
rect 2555 1579 2605 1663
rect 2641 2160 2691 2285
rect 2641 2126 2649 2160
rect 2683 2126 2691 2160
rect 2641 2092 2691 2126
rect 2641 2058 2649 2092
rect 2683 2058 2691 2092
rect 2641 2024 2691 2058
rect 2641 1990 2649 2024
rect 2683 1990 2691 2024
rect 2641 1613 2691 1990
rect 2641 1579 2649 1613
rect 2683 1579 2691 1613
rect 2727 2160 2777 2285
rect 2727 2126 2735 2160
rect 2769 2126 2777 2160
rect 2727 2092 2777 2126
rect 2727 2058 2735 2092
rect 2769 2058 2777 2092
rect 2727 2024 2777 2058
rect 2727 1990 2735 2024
rect 2769 1990 2777 2024
rect 2727 1697 2777 1990
rect 2727 1663 2735 1697
rect 2769 1663 2777 1697
rect 2727 1579 2777 1663
rect 2813 2160 2863 2285
rect 2813 2126 2821 2160
rect 2855 2126 2863 2160
rect 2813 2092 2863 2126
rect 2813 2058 2821 2092
rect 2855 2058 2863 2092
rect 2813 2024 2863 2058
rect 2813 1990 2821 2024
rect 2855 1990 2863 2024
rect 2813 1613 2863 1990
rect 2813 1579 2821 1613
rect 2855 1579 2863 1613
rect 2899 2160 2949 2285
rect 2899 2126 2907 2160
rect 2941 2126 2949 2160
rect 2899 2092 2949 2126
rect 2899 2058 2907 2092
rect 2941 2058 2949 2092
rect 2899 2024 2949 2058
rect 2899 1990 2907 2024
rect 2941 1990 2949 2024
rect 2899 1697 2949 1990
rect 2899 1663 2907 1697
rect 2941 1663 2949 1697
rect 2899 1579 2949 1663
rect 2985 2160 3035 2285
rect 2985 2126 2993 2160
rect 3027 2126 3035 2160
rect 2985 2092 3035 2126
rect 2985 2058 2993 2092
rect 3027 2058 3035 2092
rect 2985 2024 3035 2058
rect 2985 1990 2993 2024
rect 3027 1990 3035 2024
rect 2985 1613 3035 1990
rect 2985 1579 2993 1613
rect 3027 1579 3035 1613
rect 3071 2160 3121 2285
rect 3071 2126 3079 2160
rect 3113 2126 3121 2160
rect 3071 2092 3121 2126
rect 3071 2058 3079 2092
rect 3113 2058 3121 2092
rect 3071 2024 3121 2058
rect 3071 1990 3079 2024
rect 3113 1990 3121 2024
rect 3071 1697 3121 1990
rect 3071 1663 3079 1697
rect 3113 1663 3121 1697
rect 3071 1579 3121 1663
rect 577 1529 627 1579
rect 577 1495 585 1529
rect 619 1495 627 1529
rect 835 1495 843 1529
rect 877 1495 885 1529
rect 319 1277 369 1445
rect 319 1243 327 1277
rect 361 1243 369 1277
rect 319 1034 369 1243
rect 319 1000 327 1034
rect 361 1000 369 1034
rect 319 966 369 1000
rect 319 932 327 966
rect 361 932 369 966
rect 319 898 369 932
rect 319 864 327 898
rect 361 864 369 898
rect 319 739 369 864
rect 405 1361 455 1445
rect 405 1327 413 1361
rect 447 1327 455 1361
rect 405 1034 455 1327
rect 405 1000 413 1034
rect 447 1000 455 1034
rect 405 966 455 1000
rect 405 932 413 966
rect 447 932 455 966
rect 405 898 455 932
rect 405 864 413 898
rect 447 864 455 898
rect 405 739 455 864
rect 491 1277 541 1445
rect 491 1243 499 1277
rect 533 1243 541 1277
rect 491 1034 541 1243
rect 491 1000 499 1034
rect 533 1000 541 1034
rect 491 966 541 1000
rect 491 932 499 966
rect 533 932 541 966
rect 491 898 541 932
rect 491 864 499 898
rect 533 864 541 898
rect 491 739 541 864
rect 577 1411 585 1445
rect 619 1411 627 1445
rect 577 1034 627 1411
rect 577 1000 585 1034
rect 619 1000 627 1034
rect 577 966 627 1000
rect 577 932 585 966
rect 619 932 627 966
rect 577 898 627 932
rect 577 864 585 898
rect 619 864 627 898
rect 577 739 627 864
rect 663 1277 713 1445
rect 835 1361 885 1495
rect 921 1445 971 1579
rect 2469 1529 2519 1579
rect 2469 1495 2477 1529
rect 2511 1495 2519 1529
rect 921 1411 929 1445
rect 963 1411 971 1445
rect 835 1327 843 1361
rect 877 1327 885 1361
rect 1007 1361 1057 1445
rect 1007 1327 1015 1361
rect 1049 1327 1057 1361
rect 663 1243 671 1277
rect 705 1243 713 1277
rect 663 1034 713 1243
rect 663 1000 671 1034
rect 705 1000 713 1034
rect 663 966 713 1000
rect 663 932 671 966
rect 705 932 713 966
rect 663 898 713 932
rect 663 864 671 898
rect 705 864 713 898
rect 663 739 713 864
rect 1007 1034 1057 1327
rect 1007 1000 1015 1034
rect 1049 1000 1057 1034
rect 1007 966 1057 1000
rect 1007 932 1015 966
rect 1049 932 1057 966
rect 1007 898 1057 932
rect 1007 864 1015 898
rect 1049 864 1057 898
rect 1007 739 1057 864
rect 1093 1411 1101 1445
rect 1135 1411 1143 1445
rect 1093 1034 1143 1411
rect 1093 1000 1101 1034
rect 1135 1000 1143 1034
rect 1093 966 1143 1000
rect 1093 932 1101 966
rect 1135 932 1143 966
rect 1093 898 1143 932
rect 1093 864 1101 898
rect 1135 864 1143 898
rect 1093 739 1143 864
rect 1179 1361 1229 1445
rect 1179 1327 1187 1361
rect 1221 1327 1229 1361
rect 1179 1034 1229 1327
rect 1179 1000 1187 1034
rect 1221 1000 1229 1034
rect 1179 966 1229 1000
rect 1179 932 1187 966
rect 1221 932 1229 966
rect 1179 898 1229 932
rect 1179 864 1187 898
rect 1221 864 1229 898
rect 1179 739 1229 864
rect 1265 1411 1273 1445
rect 1307 1411 1315 1445
rect 1265 1034 1315 1411
rect 1265 1000 1273 1034
rect 1307 1000 1315 1034
rect 1265 966 1315 1000
rect 1265 932 1273 966
rect 1307 932 1315 966
rect 1265 898 1315 932
rect 1265 864 1273 898
rect 1307 864 1315 898
rect 1265 739 1315 864
rect 1351 1361 1401 1445
rect 1351 1327 1359 1361
rect 1393 1327 1401 1361
rect 1351 1034 1401 1327
rect 1351 1000 1359 1034
rect 1393 1000 1401 1034
rect 1351 966 1401 1000
rect 1351 932 1359 966
rect 1393 932 1401 966
rect 1351 898 1401 932
rect 1351 864 1359 898
rect 1393 864 1401 898
rect 1351 739 1401 864
rect 1437 1411 1445 1445
rect 1479 1411 1487 1445
rect 1437 1034 1487 1411
rect 1437 1000 1445 1034
rect 1479 1000 1487 1034
rect 1437 966 1487 1000
rect 1437 932 1445 966
rect 1479 932 1487 966
rect 1437 898 1487 932
rect 1437 864 1445 898
rect 1479 864 1487 898
rect 1437 739 1487 864
rect 1523 1361 1573 1445
rect 1523 1327 1531 1361
rect 1565 1327 1573 1361
rect 1523 1034 1573 1327
rect 1523 1000 1531 1034
rect 1565 1000 1573 1034
rect 1523 966 1573 1000
rect 1523 932 1531 966
rect 1565 932 1573 966
rect 1523 898 1573 932
rect 1523 864 1531 898
rect 1565 864 1573 898
rect 1523 739 1573 864
rect 1609 1411 1617 1445
rect 1651 1411 1659 1445
rect 1609 1034 1659 1411
rect 1609 1000 1617 1034
rect 1651 1000 1659 1034
rect 1609 966 1659 1000
rect 1609 932 1617 966
rect 1651 932 1659 966
rect 1609 898 1659 932
rect 1609 864 1617 898
rect 1651 864 1659 898
rect 1609 739 1659 864
rect 1695 1361 1745 1445
rect 1695 1327 1703 1361
rect 1737 1327 1745 1361
rect 1695 1034 1745 1327
rect 1695 1000 1703 1034
rect 1737 1000 1745 1034
rect 1695 966 1745 1000
rect 1695 932 1703 966
rect 1737 932 1745 966
rect 1695 898 1745 932
rect 1695 864 1703 898
rect 1737 864 1745 898
rect 1695 739 1745 864
rect 1781 1411 1789 1445
rect 1823 1411 1831 1445
rect 1781 1034 1831 1411
rect 1781 1000 1789 1034
rect 1823 1000 1831 1034
rect 1781 966 1831 1000
rect 1781 932 1789 966
rect 1823 932 1831 966
rect 1781 898 1831 932
rect 1781 864 1789 898
rect 1823 864 1831 898
rect 1781 739 1831 864
rect 1867 1361 1917 1445
rect 1867 1327 1875 1361
rect 1909 1327 1917 1361
rect 1867 1034 1917 1327
rect 1867 1000 1875 1034
rect 1909 1000 1917 1034
rect 1867 966 1917 1000
rect 1867 932 1875 966
rect 1909 932 1917 966
rect 1867 898 1917 932
rect 1867 864 1875 898
rect 1909 864 1917 898
rect 1867 739 1917 864
rect 1953 1411 1961 1445
rect 1995 1411 2003 1445
rect 1953 1034 2003 1411
rect 1953 1000 1961 1034
rect 1995 1000 2003 1034
rect 1953 966 2003 1000
rect 1953 932 1961 966
rect 1995 932 2003 966
rect 1953 898 2003 932
rect 1953 864 1961 898
rect 1995 864 2003 898
rect 1953 739 2003 864
rect 2039 1361 2089 1445
rect 2039 1327 2047 1361
rect 2081 1327 2089 1361
rect 2039 1034 2089 1327
rect 2039 1000 2047 1034
rect 2081 1000 2089 1034
rect 2039 966 2089 1000
rect 2039 932 2047 966
rect 2081 932 2089 966
rect 2039 898 2089 932
rect 2039 864 2047 898
rect 2081 864 2089 898
rect 2039 739 2089 864
rect 2383 1277 2433 1445
rect 2383 1243 2391 1277
rect 2425 1243 2433 1277
rect 2383 1034 2433 1243
rect 2383 1000 2391 1034
rect 2425 1000 2433 1034
rect 2383 966 2433 1000
rect 2383 932 2391 966
rect 2425 932 2433 966
rect 2383 898 2433 932
rect 2383 864 2391 898
rect 2425 864 2433 898
rect 2383 739 2433 864
rect 2469 1361 2519 1445
rect 2469 1327 2477 1361
rect 2511 1327 2519 1361
rect 2469 1034 2519 1327
rect 2469 1000 2477 1034
rect 2511 1000 2519 1034
rect 2469 966 2519 1000
rect 2469 932 2477 966
rect 2511 932 2519 966
rect 2469 898 2519 932
rect 2469 864 2477 898
rect 2511 864 2519 898
rect 2469 739 2519 864
rect 2555 1277 2605 1445
rect 2555 1243 2563 1277
rect 2597 1243 2605 1277
rect 2555 1034 2605 1243
rect 2555 1000 2563 1034
rect 2597 1000 2605 1034
rect 2555 966 2605 1000
rect 2555 932 2563 966
rect 2597 932 2605 966
rect 2555 898 2605 932
rect 2555 864 2563 898
rect 2597 864 2605 898
rect 2555 739 2605 864
rect 2641 1411 2649 1445
rect 2683 1411 2691 1445
rect 2641 1034 2691 1411
rect 2641 1000 2649 1034
rect 2683 1000 2691 1034
rect 2641 966 2691 1000
rect 2641 932 2649 966
rect 2683 932 2691 966
rect 2641 898 2691 932
rect 2641 864 2649 898
rect 2683 864 2691 898
rect 2641 739 2691 864
rect 2727 1277 2777 1445
rect 2727 1243 2735 1277
rect 2769 1243 2777 1277
rect 2727 1034 2777 1243
rect 2727 1000 2735 1034
rect 2769 1000 2777 1034
rect 2727 966 2777 1000
rect 2727 932 2735 966
rect 2769 932 2777 966
rect 2727 898 2777 932
rect 2727 864 2735 898
rect 2769 864 2777 898
rect 2727 739 2777 864
rect 2813 1411 2821 1445
rect 2855 1411 2863 1445
rect 2813 1034 2863 1411
rect 2813 1000 2821 1034
rect 2855 1000 2863 1034
rect 2813 966 2863 1000
rect 2813 932 2821 966
rect 2855 932 2863 966
rect 2813 898 2863 932
rect 2813 864 2821 898
rect 2855 864 2863 898
rect 2813 739 2863 864
rect 2899 1277 2949 1445
rect 2899 1243 2907 1277
rect 2941 1243 2949 1277
rect 2899 1034 2949 1243
rect 2899 1000 2907 1034
rect 2941 1000 2949 1034
rect 2899 966 2949 1000
rect 2899 932 2907 966
rect 2941 932 2949 966
rect 2899 898 2949 932
rect 2899 864 2907 898
rect 2941 864 2949 898
rect 2899 739 2949 864
rect 2985 1361 3035 1445
rect 2985 1327 2993 1361
rect 3027 1327 3035 1361
rect 2985 1034 3035 1327
rect 2985 1000 2993 1034
rect 3027 1000 3035 1034
rect 2985 966 3035 1000
rect 2985 932 2993 966
rect 3027 932 3035 966
rect 2985 898 3035 932
rect 2985 864 2993 898
rect 3027 864 3035 898
rect 2985 739 3035 864
rect 3071 1277 3121 1445
rect 3071 1243 3079 1277
rect 3113 1243 3121 1277
rect 3071 1034 3121 1243
rect 3071 1000 3079 1034
rect 3113 1000 3121 1034
rect 3071 966 3121 1000
rect 3071 932 3079 966
rect 3113 932 3121 966
rect 3071 898 3121 932
rect 3071 864 3079 898
rect 3113 864 3121 898
rect 3071 739 3121 864
rect 405 605 455 689
rect 405 571 413 605
rect 447 571 455 605
rect 405 487 455 571
rect 577 605 627 689
rect 577 571 585 605
rect 619 571 627 605
rect 577 487 627 571
rect 1093 605 1143 689
rect 1093 571 1101 605
rect 1135 571 1143 605
rect 1093 487 1143 571
rect 1265 605 1315 689
rect 1265 571 1273 605
rect 1307 571 1315 605
rect 1265 487 1315 571
rect 1437 605 1487 689
rect 1437 571 1445 605
rect 1479 571 1487 605
rect 1437 487 1487 571
rect 1609 605 1659 689
rect 1609 571 1617 605
rect 1651 571 1659 605
rect 1609 487 1659 571
rect 1781 605 1831 689
rect 1781 571 1789 605
rect 1823 571 1831 605
rect 1781 487 1831 571
rect 1953 605 2003 689
rect 1953 571 1961 605
rect 1995 571 2003 605
rect 1953 487 2003 571
rect 2469 605 2519 689
rect 2469 571 2477 605
rect 2511 571 2519 605
rect 2469 487 2519 571
rect 2641 605 2691 689
rect 2641 571 2649 605
rect 2683 571 2691 605
rect 2641 487 2691 571
rect 2813 605 2863 689
rect 2813 571 2821 605
rect 2855 571 2863 605
rect 2813 487 2863 571
rect 2985 605 3035 689
rect 2985 571 2993 605
rect 3027 571 3035 605
rect 2985 487 3035 571
rect 405 185 455 269
rect 405 151 413 185
rect 447 151 455 185
rect 405 67 455 151
rect 577 185 627 269
rect 577 151 585 185
rect 619 151 627 185
rect 577 67 627 151
rect 1093 185 1143 269
rect 1093 151 1101 185
rect 1135 151 1143 185
rect 1093 67 1143 151
rect 1265 185 1315 269
rect 1265 151 1273 185
rect 1307 151 1315 185
rect 1265 67 1315 151
rect 1437 185 1487 269
rect 1437 151 1445 185
rect 1479 151 1487 185
rect 1437 67 1487 151
rect 1609 185 1659 269
rect 1609 151 1617 185
rect 1651 151 1659 185
rect 1609 67 1659 151
rect 1781 185 1831 269
rect 1781 151 1789 185
rect 1823 151 1831 185
rect 1781 67 1831 151
rect 1953 185 2003 269
rect 1953 151 1961 185
rect 1995 151 2003 185
rect 1953 67 2003 151
rect 2469 185 2519 269
rect 2469 151 2477 185
rect 2511 151 2519 185
rect 2469 67 2519 151
rect 2641 185 2691 269
rect 2641 151 2649 185
rect 2683 151 2691 185
rect 2641 67 2691 151
rect 2813 185 2863 269
rect 2813 151 2821 185
rect 2855 151 2863 185
rect 2813 67 2863 151
rect 2985 185 3035 269
rect 2985 151 2993 185
rect 3027 151 3035 185
rect 2985 67 3035 151
<< viali >>
rect 241 2839 275 2873
rect 413 2839 447 2873
rect 413 2755 447 2789
rect 757 2839 791 2873
rect 1273 2839 1307 2873
rect 1789 2839 1823 2873
rect 1961 2839 1995 2873
rect 2133 2839 2167 2873
rect 2649 2839 2683 2873
rect 2821 2839 2855 2873
rect 2993 2839 3027 2873
rect 241 2419 275 2453
rect 757 2419 791 2453
rect 1273 2419 1307 2453
rect 1703 2419 1737 2453
rect 1703 2335 1737 2369
rect 1789 2419 1823 2453
rect 1961 2419 1995 2453
rect 2133 2419 2167 2453
rect 2649 2419 2683 2453
rect 2821 2419 2855 2453
rect 2993 2419 3027 2453
rect 155 1663 189 1697
rect 241 1579 275 1613
rect 327 1663 361 1697
rect 671 1663 705 1697
rect 585 1579 619 1613
rect 757 1579 791 1613
rect 843 1663 877 1697
rect 1187 1663 1221 1697
rect 929 1579 963 1613
rect 1273 1579 1307 1613
rect 1359 1663 1393 1697
rect 1703 1663 1737 1697
rect 1789 1579 1823 1613
rect 1875 1663 1909 1697
rect 1961 1579 1995 1613
rect 2047 1663 2081 1697
rect 2133 1579 2167 1613
rect 2219 1663 2253 1697
rect 2563 1663 2597 1697
rect 2477 1579 2511 1613
rect 2649 1579 2683 1613
rect 2735 1663 2769 1697
rect 2821 1579 2855 1613
rect 2907 1663 2941 1697
rect 2993 1579 3027 1613
rect 3079 1663 3113 1697
rect 585 1495 619 1529
rect 843 1495 877 1529
rect 327 1243 361 1277
rect 413 1327 447 1361
rect 499 1243 533 1277
rect 585 1411 619 1445
rect 2477 1495 2511 1529
rect 929 1411 963 1445
rect 843 1327 877 1361
rect 1015 1327 1049 1361
rect 671 1243 705 1277
rect 1101 1411 1135 1445
rect 1187 1327 1221 1361
rect 1273 1411 1307 1445
rect 1359 1327 1393 1361
rect 1445 1411 1479 1445
rect 1531 1327 1565 1361
rect 1617 1411 1651 1445
rect 1703 1327 1737 1361
rect 1789 1411 1823 1445
rect 1875 1327 1909 1361
rect 1961 1411 1995 1445
rect 2047 1327 2081 1361
rect 2391 1243 2425 1277
rect 2477 1327 2511 1361
rect 2563 1243 2597 1277
rect 2649 1411 2683 1445
rect 2735 1243 2769 1277
rect 2821 1411 2855 1445
rect 2907 1243 2941 1277
rect 2993 1327 3027 1361
rect 3079 1243 3113 1277
rect 413 571 447 605
rect 585 571 619 605
rect 1101 571 1135 605
rect 1273 571 1307 605
rect 1445 571 1479 605
rect 1617 571 1651 605
rect 1789 571 1823 605
rect 1961 571 1995 605
rect 2477 571 2511 605
rect 2649 571 2683 605
rect 2821 571 2855 605
rect 2993 571 3027 605
rect 413 151 447 185
rect 585 151 619 185
rect 1101 151 1135 185
rect 1273 151 1307 185
rect 1445 151 1479 185
rect 1617 151 1651 185
rect 1789 151 1823 185
rect 1961 151 1995 185
rect 2477 151 2511 185
rect 2649 151 2683 185
rect 2821 151 2855 185
rect 2993 151 3027 185
<< metal1 >>
rect 224 2873 464 2884
rect 224 2839 241 2873
rect 275 2839 413 2873
rect 447 2839 464 2873
rect 224 2828 464 2839
rect 654 2882 894 2884
rect 654 2873 834 2882
rect 654 2839 757 2873
rect 791 2839 834 2873
rect 654 2830 834 2839
rect 886 2830 894 2882
rect 654 2828 894 2830
rect 1170 2882 1410 2884
rect 1170 2830 1178 2882
rect 1230 2873 1410 2882
rect 1230 2839 1273 2873
rect 1307 2839 1410 2873
rect 1230 2830 1410 2839
rect 1170 2828 1410 2830
rect 1602 2882 3044 2884
rect 1602 2830 1608 2882
rect 1660 2873 3044 2882
rect 1660 2839 1789 2873
rect 1823 2839 1961 2873
rect 1995 2839 2133 2873
rect 2167 2839 2649 2873
rect 2683 2839 2821 2873
rect 2855 2839 2993 2873
rect 3027 2839 3044 2873
rect 1660 2830 3044 2839
rect 1602 2828 3044 2830
rect 396 2798 892 2800
rect 396 2789 834 2798
rect 396 2755 413 2789
rect 447 2755 834 2789
rect 396 2746 834 2755
rect 886 2746 892 2798
rect 396 2744 892 2746
rect 224 2462 808 2464
rect 224 2453 318 2462
rect 224 2419 241 2453
rect 275 2419 318 2453
rect 224 2410 318 2419
rect 370 2453 808 2462
rect 370 2419 757 2453
rect 791 2419 808 2453
rect 370 2410 808 2419
rect 224 2408 808 2410
rect 1256 2462 1496 2464
rect 1256 2410 1264 2462
rect 1316 2410 1496 2462
rect 1256 2408 1496 2410
rect 1686 2453 2184 2464
rect 1686 2419 1703 2453
rect 1737 2419 1789 2453
rect 1823 2419 1961 2453
rect 1995 2419 2133 2453
rect 2167 2419 2184 2453
rect 1686 2408 2184 2419
rect 2632 2453 3044 2464
rect 2632 2419 2649 2453
rect 2683 2419 2821 2453
rect 2855 2419 2993 2453
rect 3027 2419 3044 2453
rect 2632 2408 3044 2419
rect 1258 2378 1754 2380
rect 1258 2326 1264 2378
rect 1316 2369 1754 2378
rect 1316 2335 1703 2369
rect 1737 2335 1754 2369
rect 1316 2326 1754 2335
rect 1258 2324 1754 2326
rect 828 1790 1236 1792
rect 828 1738 834 1790
rect 886 1738 1178 1790
rect 1230 1738 1236 1790
rect 828 1736 1236 1738
rect 138 1706 378 1708
rect 138 1697 232 1706
rect 138 1663 155 1697
rect 189 1663 232 1697
rect 138 1654 232 1663
rect 284 1697 378 1706
rect 284 1663 327 1697
rect 361 1663 378 1697
rect 284 1654 378 1663
rect 138 1652 378 1654
rect 654 1706 894 1708
rect 654 1697 834 1706
rect 654 1663 671 1697
rect 705 1663 834 1697
rect 654 1654 834 1663
rect 886 1654 894 1706
rect 654 1652 894 1654
rect 1170 1706 1410 1708
rect 1170 1654 1178 1706
rect 1230 1697 1410 1706
rect 1230 1663 1359 1697
rect 1393 1663 1410 1697
rect 1230 1654 1410 1663
rect 1170 1652 1410 1654
rect 1686 1706 3130 1708
rect 1686 1697 2468 1706
rect 1686 1663 1703 1697
rect 1737 1663 1875 1697
rect 1909 1663 2047 1697
rect 2081 1663 2219 1697
rect 2253 1663 2468 1697
rect 1686 1654 2468 1663
rect 2520 1697 3130 1706
rect 2520 1663 2563 1697
rect 2597 1663 2735 1697
rect 2769 1663 2907 1697
rect 2941 1663 3079 1697
rect 3113 1663 3130 1697
rect 2520 1654 3130 1663
rect 1686 1652 3130 1654
rect 224 1622 464 1624
rect 224 1570 232 1622
rect 284 1570 464 1622
rect 224 1568 464 1570
rect 568 1613 980 1624
rect 568 1579 585 1613
rect 619 1579 757 1613
rect 791 1579 929 1613
rect 963 1579 980 1613
rect 568 1568 980 1579
rect 1256 1622 1496 1624
rect 1256 1570 1264 1622
rect 1316 1570 1496 1622
rect 1256 1568 1496 1570
rect 1688 1622 2184 1624
rect 1688 1570 1694 1622
rect 1746 1613 2184 1622
rect 1746 1579 1789 1613
rect 1823 1579 1961 1613
rect 1995 1579 2133 1613
rect 2167 1579 2184 1613
rect 1746 1570 2184 1579
rect 1688 1568 2184 1570
rect 2460 1613 3044 1624
rect 2460 1579 2477 1613
rect 2511 1579 2649 1613
rect 2683 1579 2821 1613
rect 2855 1579 2993 1613
rect 3027 1579 3044 1613
rect 2460 1568 3044 1579
rect 226 1538 636 1540
rect 226 1486 232 1538
rect 284 1529 636 1538
rect 284 1495 585 1529
rect 619 1495 636 1529
rect 284 1486 636 1495
rect 226 1484 636 1486
rect 826 1529 2528 1540
rect 826 1495 843 1529
rect 877 1495 2477 1529
rect 2511 1495 2528 1529
rect 826 1484 2528 1495
rect 568 1454 808 1456
rect 568 1402 576 1454
rect 628 1402 808 1454
rect 568 1400 808 1402
rect 912 1445 2012 1456
rect 912 1411 929 1445
rect 963 1411 1101 1445
rect 1135 1411 1273 1445
rect 1307 1411 1445 1445
rect 1479 1411 1617 1445
rect 1651 1411 1789 1445
rect 1823 1411 1961 1445
rect 1995 1411 2012 1445
rect 912 1400 2012 1411
rect 2632 1454 2872 1456
rect 2632 1402 2640 1454
rect 2692 1445 2872 1454
rect 2692 1411 2821 1445
rect 2855 1411 2872 1445
rect 2692 1402 2872 1411
rect 2632 1400 2872 1402
rect 312 1370 894 1372
rect 312 1318 318 1370
rect 370 1361 894 1370
rect 370 1327 413 1361
rect 447 1327 843 1361
rect 877 1327 894 1361
rect 370 1318 894 1327
rect 312 1316 894 1318
rect 998 1370 2098 1372
rect 998 1361 1608 1370
rect 998 1327 1015 1361
rect 1049 1327 1187 1361
rect 1221 1327 1359 1361
rect 1393 1327 1531 1361
rect 1565 1327 1608 1361
rect 998 1318 1608 1327
rect 1660 1361 2098 1370
rect 1660 1327 1703 1361
rect 1737 1327 1875 1361
rect 1909 1327 2047 1361
rect 2081 1327 2098 1361
rect 1660 1318 2098 1327
rect 998 1316 2098 1318
rect 2460 1370 3044 1372
rect 2460 1318 2468 1370
rect 2520 1361 3044 1370
rect 2520 1327 2993 1361
rect 3027 1327 3044 1361
rect 2520 1318 3044 1327
rect 2460 1316 3044 1318
rect 310 1286 722 1288
rect 310 1277 404 1286
rect 310 1243 327 1277
rect 361 1243 404 1277
rect 310 1234 404 1243
rect 456 1277 722 1286
rect 456 1243 499 1277
rect 533 1243 671 1277
rect 705 1243 722 1277
rect 456 1234 722 1243
rect 310 1232 722 1234
rect 2374 1286 3130 1288
rect 2374 1277 2812 1286
rect 2374 1243 2391 1277
rect 2425 1243 2563 1277
rect 2597 1243 2735 1277
rect 2769 1243 2812 1277
rect 2374 1234 2812 1243
rect 2864 1277 3130 1286
rect 2864 1243 2907 1277
rect 2941 1243 3079 1277
rect 3113 1243 3130 1277
rect 2864 1234 3130 1243
rect 2374 1232 3130 1234
rect 2290 698 2698 700
rect 2290 646 2296 698
rect 2348 646 2640 698
rect 2692 646 2698 698
rect 2290 644 2698 646
rect 396 614 636 616
rect 396 605 576 614
rect 396 571 413 605
rect 447 571 576 605
rect 396 562 576 571
rect 628 562 636 614
rect 396 560 636 562
rect 1084 614 2354 616
rect 1084 605 1264 614
rect 1316 605 2296 614
rect 1084 571 1101 605
rect 1135 571 1264 605
rect 1316 571 1445 605
rect 1479 571 1617 605
rect 1651 571 1789 605
rect 1823 571 1961 605
rect 1995 571 2296 605
rect 1084 562 1264 571
rect 1316 562 2296 571
rect 2348 562 2354 614
rect 1084 560 2354 562
rect 2460 614 3044 616
rect 2460 605 2640 614
rect 2692 605 3044 614
rect 2460 571 2477 605
rect 2511 571 2640 605
rect 2692 571 2821 605
rect 2855 571 2993 605
rect 3027 571 3044 605
rect 2460 562 2640 571
rect 2692 562 3044 571
rect 2460 560 3044 562
rect 1602 278 2870 280
rect 1602 226 1608 278
rect 1660 226 2812 278
rect 2864 226 2870 278
rect 1602 224 2870 226
rect 396 194 636 196
rect 396 142 404 194
rect 456 185 636 194
rect 456 151 585 185
rect 619 151 636 185
rect 456 142 636 151
rect 396 140 636 142
rect 1084 194 2012 196
rect 1084 185 1608 194
rect 1660 185 2012 194
rect 1084 151 1101 185
rect 1135 151 1273 185
rect 1307 151 1445 185
rect 1479 151 1608 185
rect 1660 151 1789 185
rect 1823 151 1961 185
rect 1995 151 2012 185
rect 1084 142 1608 151
rect 1660 142 2012 151
rect 1084 140 2012 142
rect 2460 194 3044 196
rect 2460 185 2812 194
rect 2864 185 3044 194
rect 2460 151 2477 185
rect 2511 151 2649 185
rect 2683 151 2812 185
rect 2864 151 2993 185
rect 3027 151 3044 185
rect 2460 142 2812 151
rect 2864 142 3044 151
rect 2460 140 3044 142
<< via1 >>
rect 834 2830 886 2882
rect 1178 2830 1230 2882
rect 1608 2830 1660 2882
rect 834 2746 886 2798
rect 318 2410 370 2462
rect 1264 2453 1316 2462
rect 1264 2419 1273 2453
rect 1273 2419 1307 2453
rect 1307 2419 1316 2453
rect 1264 2410 1316 2419
rect 1264 2326 1316 2378
rect 834 1738 886 1790
rect 1178 1738 1230 1790
rect 232 1654 284 1706
rect 834 1697 886 1706
rect 834 1663 843 1697
rect 843 1663 877 1697
rect 877 1663 886 1697
rect 834 1654 886 1663
rect 1178 1697 1230 1706
rect 1178 1663 1187 1697
rect 1187 1663 1221 1697
rect 1221 1663 1230 1697
rect 1178 1654 1230 1663
rect 2468 1654 2520 1706
rect 232 1613 284 1622
rect 232 1579 241 1613
rect 241 1579 275 1613
rect 275 1579 284 1613
rect 232 1570 284 1579
rect 1264 1613 1316 1622
rect 1264 1579 1273 1613
rect 1273 1579 1307 1613
rect 1307 1579 1316 1613
rect 1264 1570 1316 1579
rect 1694 1570 1746 1622
rect 232 1486 284 1538
rect 576 1445 628 1454
rect 576 1411 585 1445
rect 585 1411 619 1445
rect 619 1411 628 1445
rect 576 1402 628 1411
rect 2640 1445 2692 1454
rect 2640 1411 2649 1445
rect 2649 1411 2683 1445
rect 2683 1411 2692 1445
rect 2640 1402 2692 1411
rect 318 1318 370 1370
rect 1608 1318 1660 1370
rect 2468 1361 2520 1370
rect 2468 1327 2477 1361
rect 2477 1327 2511 1361
rect 2511 1327 2520 1361
rect 2468 1318 2520 1327
rect 404 1234 456 1286
rect 2812 1234 2864 1286
rect 2296 646 2348 698
rect 2640 646 2692 698
rect 576 605 628 614
rect 576 571 585 605
rect 585 571 619 605
rect 619 571 628 605
rect 576 562 628 571
rect 1264 605 1316 614
rect 1264 571 1273 605
rect 1273 571 1307 605
rect 1307 571 1316 605
rect 1264 562 1316 571
rect 2296 562 2348 614
rect 2640 605 2692 614
rect 2640 571 2649 605
rect 2649 571 2683 605
rect 2683 571 2692 605
rect 2640 562 2692 571
rect 1608 226 1660 278
rect 2812 226 2864 278
rect 404 185 456 194
rect 404 151 413 185
rect 413 151 447 185
rect 447 151 456 185
rect 404 142 456 151
rect 1608 185 1660 194
rect 1608 151 1617 185
rect 1617 151 1651 185
rect 1651 151 1660 185
rect 1608 142 1660 151
rect 2812 185 2864 194
rect 2812 151 2821 185
rect 2821 151 2855 185
rect 2855 151 2864 185
rect 2812 142 2864 151
<< metal2 >>
rect 832 2882 888 2888
rect 832 2830 834 2882
rect 886 2830 888 2882
rect 832 2798 888 2830
rect 832 2746 834 2798
rect 886 2746 888 2798
rect 316 2462 372 2468
rect 316 2410 318 2462
rect 370 2410 372 2462
rect 230 1706 286 1796
rect 230 1654 232 1706
rect 284 1654 286 1706
rect 230 1622 286 1654
rect 230 1570 232 1622
rect 284 1570 286 1622
rect 230 1538 286 1570
rect 230 1486 232 1538
rect 284 1486 286 1538
rect 230 1480 286 1486
rect 316 1370 372 2410
rect 832 1790 888 2746
rect 832 1738 834 1790
rect 886 1738 888 1790
rect 832 1706 888 1738
rect 832 1654 834 1706
rect 886 1654 888 1706
rect 316 1318 318 1370
rect 370 1318 372 1370
rect 316 1312 372 1318
rect 574 1540 630 1549
rect 574 1454 630 1484
rect 574 1402 576 1454
rect 628 1402 630 1454
rect 402 1288 458 1297
rect 402 194 458 1232
rect 574 614 630 1402
rect 832 1288 888 1654
rect 1176 2882 1232 2888
rect 1176 2830 1178 2882
rect 1230 2830 1232 2882
rect 1176 1790 1232 2830
rect 1606 2882 1662 2888
rect 1606 2830 1608 2882
rect 1660 2830 1662 2882
rect 1176 1738 1178 1790
rect 1230 1738 1232 1790
rect 1176 1706 1232 1738
rect 1176 1654 1178 1706
rect 1230 1654 1232 1706
rect 1176 1648 1232 1654
rect 1262 2462 1318 2468
rect 1262 2410 1264 2462
rect 1316 2410 1318 2462
rect 1262 2378 1318 2410
rect 1262 2326 1264 2378
rect 1316 2326 1318 2378
rect 832 1223 888 1232
rect 1262 1622 1318 2326
rect 1262 1570 1264 1622
rect 1316 1570 1318 1622
rect 574 562 576 614
rect 628 562 630 614
rect 574 556 630 562
rect 1262 614 1318 1570
rect 1262 562 1264 614
rect 1316 562 1318 614
rect 1262 556 1318 562
rect 1606 1370 1662 2830
rect 2466 1706 2522 1712
rect 2466 1654 2468 1706
rect 2520 1654 2522 1706
rect 1692 1622 1748 1628
rect 1692 1570 1694 1622
rect 1746 1570 1748 1622
rect 1692 1540 1748 1570
rect 1692 1475 1748 1484
rect 1606 1318 1608 1370
rect 1660 1318 1662 1370
rect 402 142 404 194
rect 456 142 458 194
rect 402 136 458 142
rect 1606 278 1662 1318
rect 2466 1370 2522 1654
rect 2466 1318 2468 1370
rect 2520 1318 2522 1370
rect 2466 1312 2522 1318
rect 2638 1454 2694 1460
rect 2638 1402 2640 1454
rect 2692 1402 2694 1454
rect 2294 698 2350 704
rect 2294 646 2296 698
rect 2348 646 2350 698
rect 2294 614 2350 646
rect 2294 562 2296 614
rect 2348 562 2350 614
rect 2294 556 2350 562
rect 2638 698 2694 1402
rect 2638 646 2640 698
rect 2692 646 2694 698
rect 2638 614 2694 646
rect 2638 562 2640 614
rect 2692 562 2694 614
rect 2638 556 2694 562
rect 2810 1286 2866 1292
rect 2810 1234 2812 1286
rect 2864 1234 2866 1286
rect 1606 226 1608 278
rect 1660 226 1662 278
rect 1606 194 1662 226
rect 1606 142 1608 194
rect 1660 142 1662 194
rect 1606 136 1662 142
rect 2810 278 2866 1234
rect 2810 226 2812 278
rect 2864 226 2866 278
rect 2810 194 2866 226
rect 2810 142 2812 194
rect 2864 142 2866 194
rect 2810 136 2866 142
<< via2 >>
rect 574 1484 630 1540
rect 402 1286 458 1288
rect 402 1234 404 1286
rect 404 1234 456 1286
rect 456 1234 458 1286
rect 402 1232 458 1234
rect 832 1232 888 1288
rect 1692 1484 1748 1540
<< metal3 >>
rect 569 1540 1753 1592
rect 569 1484 574 1540
rect 630 1484 1692 1540
rect 1748 1484 1753 1540
rect 569 1432 1753 1484
rect 397 1288 893 1340
rect 397 1232 402 1288
rect 458 1232 832 1288
rect 888 1232 893 1288
rect 397 1180 893 1232
<< labels >>
flabel locali 1093 1034 1143 1411 0 FreeSans 1600 0 0 0 vout
port 0 nsew
flabel poly 2694 2184 2724 2463 0 FreeSans 1600 0 0 0 vpos
port 1 nsew
flabel pwell 1247 2718 1333 2994 0 FreeSans 1600 0 0 0 gnd
port 2 nsew
flabel nwell 1548 0 3268 3024 0 FreeSans 1600 0 0 0 vdd
port 4 nsew
<< end >>
