magic
tech sky130A
magscale 1 2
timestamp 1678494626
<< nwell >>
rect 0 1932 3784 2688
rect 0 420 6020 1932
rect 6536 1176 11524 2688
rect 0 0 3784 420
rect 7052 0 11524 1176
<< pwell >>
rect 1161 3894 1247 4170
rect 3053 3894 3139 4170
rect 6751 3894 6837 4170
rect 9245 3894 9331 4170
rect 6235 3558 6321 3834
rect 1067 3124 1341 3386
rect 2959 3124 3233 3386
rect 4429 3138 4515 3414
rect 5547 3138 5633 3414
rect 6657 3124 6931 3386
rect 9151 3124 9425 3386
rect 6141 2788 6415 3050
rect 4335 2368 4609 2630
rect 5453 2368 5727 2630
rect 6235 2046 6321 2322
rect 6141 1276 6415 1538
<< nmos >>
rect 1146 3150 1176 3360
rect 1232 3150 1262 3360
rect 3038 3150 3068 3360
rect 3124 3150 3154 3360
rect 6736 3150 6766 3360
rect 6822 3150 6852 3360
rect 9230 3150 9260 3360
rect 9316 3150 9346 3360
rect 6220 2814 6250 3024
rect 6306 2814 6336 3024
rect 4414 2394 4444 2604
rect 4500 2394 4530 2604
rect 5532 2394 5562 2604
rect 5618 2394 5648 2604
rect 6220 1302 6250 1512
rect 6306 1302 6336 1512
<< pmos >>
rect 200 2016 230 2226
rect 286 2016 316 2226
rect 372 2016 402 2226
rect 458 2016 488 2226
rect 544 2016 574 2226
rect 630 2016 660 2226
rect 716 2016 746 2226
rect 802 2016 832 2226
rect 888 2016 918 2226
rect 974 2016 1004 2226
rect 1060 2016 1090 2226
rect 1146 2016 1176 2226
rect 1232 2016 1262 2226
rect 1318 2016 1348 2226
rect 1404 2016 1434 2226
rect 1490 2016 1520 2226
rect 1576 2016 1606 2226
rect 1662 2016 1692 2226
rect 1748 2016 1778 2226
rect 1834 2016 1864 2226
rect 1920 2016 1950 2226
rect 2006 2016 2036 2226
rect 2092 2016 2122 2226
rect 2178 2016 2208 2226
rect 2608 2016 2638 2226
rect 2694 2016 2724 2226
rect 2780 2016 2810 2226
rect 2866 2016 2896 2226
rect 2952 2016 2982 2226
rect 3038 2016 3068 2226
rect 3124 2016 3154 2226
rect 3210 2016 3240 2226
rect 3296 2016 3326 2226
rect 3382 2016 3412 2226
rect 3468 2016 3498 2226
rect 3554 2016 3584 2226
rect 6736 2016 6766 2226
rect 6822 2016 6852 2226
rect 7252 2016 7282 2226
rect 7338 2016 7368 2226
rect 7424 2016 7454 2226
rect 7510 2016 7540 2226
rect 7596 2016 7626 2226
rect 7682 2016 7712 2226
rect 7768 2016 7798 2226
rect 7854 2016 7884 2226
rect 7940 2016 7970 2226
rect 8026 2016 8056 2226
rect 8112 2016 8142 2226
rect 8198 2016 8228 2226
rect 8284 2016 8314 2226
rect 8370 2016 8400 2226
rect 8456 2016 8486 2226
rect 8542 2016 8572 2226
rect 8628 2016 8658 2226
rect 8714 2016 8744 2226
rect 8800 2016 8830 2226
rect 8886 2016 8916 2226
rect 8972 2016 9002 2226
rect 9058 2016 9088 2226
rect 9144 2016 9174 2226
rect 9230 2016 9260 2226
rect 9316 2016 9346 2226
rect 9402 2016 9432 2226
rect 9488 2016 9518 2226
rect 9574 2016 9604 2226
rect 9660 2016 9690 2226
rect 9746 2016 9776 2226
rect 9832 2016 9862 2226
rect 9918 2016 9948 2226
rect 10004 2016 10034 2226
rect 10090 2016 10120 2226
rect 10176 2016 10206 2226
rect 10262 2016 10292 2226
rect 10348 2016 10378 2226
rect 10434 2016 10464 2226
rect 10520 2016 10550 2226
rect 10606 2016 10636 2226
rect 10692 2016 10722 2226
rect 10778 2016 10808 2226
rect 10864 2016 10894 2226
rect 10950 2016 10980 2226
rect 11036 2016 11066 2226
rect 11122 2016 11152 2226
rect 11208 2016 11238 2226
rect 11294 2016 11324 2226
rect 3984 1260 4014 1470
rect 4070 1260 4100 1470
rect 4156 1260 4186 1470
rect 4242 1260 4272 1470
rect 4328 1260 4358 1470
rect 4414 1260 4444 1470
rect 4500 1260 4530 1470
rect 4586 1260 4616 1470
rect 4672 1260 4702 1470
rect 4758 1260 4788 1470
rect 4844 1260 4874 1470
rect 4930 1260 4960 1470
rect 5360 1260 5390 1470
rect 5446 1260 5476 1470
rect 5532 1260 5562 1470
rect 5618 1260 5648 1470
rect 5704 1260 5734 1470
rect 5790 1260 5820 1470
rect 200 840 230 1050
rect 286 840 316 1050
rect 372 840 402 1050
rect 458 840 488 1050
rect 544 840 574 1050
rect 630 840 660 1050
rect 716 840 746 1050
rect 802 840 832 1050
rect 888 840 918 1050
rect 974 840 1004 1050
rect 1060 840 1090 1050
rect 1146 840 1176 1050
rect 1232 840 1262 1050
rect 1318 840 1348 1050
rect 1404 840 1434 1050
rect 1490 840 1520 1050
rect 1576 840 1606 1050
rect 1662 840 1692 1050
rect 1748 840 1778 1050
rect 1834 840 1864 1050
rect 1920 840 1950 1050
rect 2006 840 2036 1050
rect 2092 840 2122 1050
rect 2178 840 2208 1050
rect 2608 840 2638 1050
rect 2694 840 2724 1050
rect 2780 840 2810 1050
rect 2866 840 2896 1050
rect 2952 840 2982 1050
rect 3038 840 3068 1050
rect 3124 840 3154 1050
rect 3210 840 3240 1050
rect 3296 840 3326 1050
rect 3382 840 3412 1050
rect 3468 840 3498 1050
rect 3554 840 3584 1050
rect 7252 840 7282 1050
rect 7338 840 7368 1050
rect 7424 840 7454 1050
rect 7510 840 7540 1050
rect 7596 840 7626 1050
rect 7682 840 7712 1050
rect 7768 840 7798 1050
rect 7854 840 7884 1050
rect 7940 840 7970 1050
rect 8026 840 8056 1050
rect 8112 840 8142 1050
rect 8198 840 8228 1050
rect 8284 840 8314 1050
rect 8370 840 8400 1050
rect 8456 840 8486 1050
rect 8542 840 8572 1050
rect 8628 840 8658 1050
rect 8714 840 8744 1050
rect 8800 840 8830 1050
rect 8886 840 8916 1050
rect 8972 840 9002 1050
rect 9058 840 9088 1050
rect 9144 840 9174 1050
rect 9230 840 9260 1050
rect 9316 840 9346 1050
rect 9402 840 9432 1050
rect 9488 840 9518 1050
rect 9574 840 9604 1050
rect 9660 840 9690 1050
rect 9746 840 9776 1050
rect 9832 840 9862 1050
rect 9918 840 9948 1050
rect 10004 840 10034 1050
rect 10090 840 10120 1050
rect 10176 840 10206 1050
rect 10262 840 10292 1050
rect 10348 840 10378 1050
rect 10434 840 10464 1050
rect 10520 840 10550 1050
rect 10606 840 10636 1050
rect 10692 840 10722 1050
rect 10778 840 10808 1050
rect 10864 840 10894 1050
rect 10950 840 10980 1050
rect 11036 840 11066 1050
rect 11122 840 11152 1050
rect 11208 840 11238 1050
rect 11294 840 11324 1050
<< ndiff >>
rect 1093 3336 1146 3360
rect 1093 3302 1101 3336
rect 1135 3302 1146 3336
rect 1093 3268 1146 3302
rect 1093 3234 1101 3268
rect 1135 3234 1146 3268
rect 1093 3200 1146 3234
rect 1093 3166 1101 3200
rect 1135 3166 1146 3200
rect 1093 3150 1146 3166
rect 1176 3336 1232 3360
rect 1176 3302 1187 3336
rect 1221 3302 1232 3336
rect 1176 3268 1232 3302
rect 1176 3234 1187 3268
rect 1221 3234 1232 3268
rect 1176 3200 1232 3234
rect 1176 3166 1187 3200
rect 1221 3166 1232 3200
rect 1176 3150 1232 3166
rect 1262 3336 1315 3360
rect 1262 3302 1273 3336
rect 1307 3302 1315 3336
rect 1262 3268 1315 3302
rect 1262 3234 1273 3268
rect 1307 3234 1315 3268
rect 1262 3200 1315 3234
rect 1262 3166 1273 3200
rect 1307 3166 1315 3200
rect 1262 3150 1315 3166
rect 2985 3336 3038 3360
rect 2985 3302 2993 3336
rect 3027 3302 3038 3336
rect 2985 3268 3038 3302
rect 2985 3234 2993 3268
rect 3027 3234 3038 3268
rect 2985 3200 3038 3234
rect 2985 3166 2993 3200
rect 3027 3166 3038 3200
rect 2985 3150 3038 3166
rect 3068 3336 3124 3360
rect 3068 3302 3079 3336
rect 3113 3302 3124 3336
rect 3068 3268 3124 3302
rect 3068 3234 3079 3268
rect 3113 3234 3124 3268
rect 3068 3200 3124 3234
rect 3068 3166 3079 3200
rect 3113 3166 3124 3200
rect 3068 3150 3124 3166
rect 3154 3336 3207 3360
rect 3154 3302 3165 3336
rect 3199 3302 3207 3336
rect 3154 3268 3207 3302
rect 3154 3234 3165 3268
rect 3199 3234 3207 3268
rect 3154 3200 3207 3234
rect 3154 3166 3165 3200
rect 3199 3166 3207 3200
rect 3154 3150 3207 3166
rect 6683 3336 6736 3360
rect 6683 3302 6691 3336
rect 6725 3302 6736 3336
rect 6683 3268 6736 3302
rect 6683 3234 6691 3268
rect 6725 3234 6736 3268
rect 6683 3200 6736 3234
rect 6683 3166 6691 3200
rect 6725 3166 6736 3200
rect 6683 3150 6736 3166
rect 6766 3336 6822 3360
rect 6766 3302 6777 3336
rect 6811 3302 6822 3336
rect 6766 3268 6822 3302
rect 6766 3234 6777 3268
rect 6811 3234 6822 3268
rect 6766 3200 6822 3234
rect 6766 3166 6777 3200
rect 6811 3166 6822 3200
rect 6766 3150 6822 3166
rect 6852 3336 6905 3360
rect 6852 3302 6863 3336
rect 6897 3302 6905 3336
rect 6852 3268 6905 3302
rect 6852 3234 6863 3268
rect 6897 3234 6905 3268
rect 6852 3200 6905 3234
rect 6852 3166 6863 3200
rect 6897 3166 6905 3200
rect 6852 3150 6905 3166
rect 9177 3336 9230 3360
rect 9177 3302 9185 3336
rect 9219 3302 9230 3336
rect 9177 3268 9230 3302
rect 9177 3234 9185 3268
rect 9219 3234 9230 3268
rect 9177 3200 9230 3234
rect 9177 3166 9185 3200
rect 9219 3166 9230 3200
rect 9177 3150 9230 3166
rect 9260 3336 9316 3360
rect 9260 3302 9271 3336
rect 9305 3302 9316 3336
rect 9260 3268 9316 3302
rect 9260 3234 9271 3268
rect 9305 3234 9316 3268
rect 9260 3200 9316 3234
rect 9260 3166 9271 3200
rect 9305 3166 9316 3200
rect 9260 3150 9316 3166
rect 9346 3336 9399 3360
rect 9346 3302 9357 3336
rect 9391 3302 9399 3336
rect 9346 3268 9399 3302
rect 9346 3234 9357 3268
rect 9391 3234 9399 3268
rect 9346 3200 9399 3234
rect 9346 3166 9357 3200
rect 9391 3166 9399 3200
rect 9346 3150 9399 3166
rect 6167 3000 6220 3024
rect 6167 2966 6175 3000
rect 6209 2966 6220 3000
rect 6167 2932 6220 2966
rect 6167 2898 6175 2932
rect 6209 2898 6220 2932
rect 6167 2864 6220 2898
rect 6167 2830 6175 2864
rect 6209 2830 6220 2864
rect 6167 2814 6220 2830
rect 6250 3000 6306 3024
rect 6250 2966 6261 3000
rect 6295 2966 6306 3000
rect 6250 2932 6306 2966
rect 6250 2898 6261 2932
rect 6295 2898 6306 2932
rect 6250 2864 6306 2898
rect 6250 2830 6261 2864
rect 6295 2830 6306 2864
rect 6250 2814 6306 2830
rect 6336 3000 6389 3024
rect 6336 2966 6347 3000
rect 6381 2966 6389 3000
rect 6336 2932 6389 2966
rect 6336 2898 6347 2932
rect 6381 2898 6389 2932
rect 6336 2864 6389 2898
rect 6336 2830 6347 2864
rect 6381 2830 6389 2864
rect 6336 2814 6389 2830
rect 4361 2580 4414 2604
rect 4361 2546 4369 2580
rect 4403 2546 4414 2580
rect 4361 2512 4414 2546
rect 4361 2478 4369 2512
rect 4403 2478 4414 2512
rect 4361 2444 4414 2478
rect 4361 2410 4369 2444
rect 4403 2410 4414 2444
rect 4361 2394 4414 2410
rect 4444 2580 4500 2604
rect 4444 2546 4455 2580
rect 4489 2546 4500 2580
rect 4444 2512 4500 2546
rect 4444 2478 4455 2512
rect 4489 2478 4500 2512
rect 4444 2444 4500 2478
rect 4444 2410 4455 2444
rect 4489 2410 4500 2444
rect 4444 2394 4500 2410
rect 4530 2580 4583 2604
rect 4530 2546 4541 2580
rect 4575 2546 4583 2580
rect 4530 2512 4583 2546
rect 4530 2478 4541 2512
rect 4575 2478 4583 2512
rect 4530 2444 4583 2478
rect 4530 2410 4541 2444
rect 4575 2410 4583 2444
rect 4530 2394 4583 2410
rect 5479 2580 5532 2604
rect 5479 2546 5487 2580
rect 5521 2546 5532 2580
rect 5479 2512 5532 2546
rect 5479 2478 5487 2512
rect 5521 2478 5532 2512
rect 5479 2444 5532 2478
rect 5479 2410 5487 2444
rect 5521 2410 5532 2444
rect 5479 2394 5532 2410
rect 5562 2580 5618 2604
rect 5562 2546 5573 2580
rect 5607 2546 5618 2580
rect 5562 2512 5618 2546
rect 5562 2478 5573 2512
rect 5607 2478 5618 2512
rect 5562 2444 5618 2478
rect 5562 2410 5573 2444
rect 5607 2410 5618 2444
rect 5562 2394 5618 2410
rect 5648 2580 5701 2604
rect 5648 2546 5659 2580
rect 5693 2546 5701 2580
rect 5648 2512 5701 2546
rect 5648 2478 5659 2512
rect 5693 2478 5701 2512
rect 5648 2444 5701 2478
rect 5648 2410 5659 2444
rect 5693 2410 5701 2444
rect 5648 2394 5701 2410
rect 6167 1488 6220 1512
rect 6167 1454 6175 1488
rect 6209 1454 6220 1488
rect 6167 1420 6220 1454
rect 6167 1386 6175 1420
rect 6209 1386 6220 1420
rect 6167 1352 6220 1386
rect 6167 1318 6175 1352
rect 6209 1318 6220 1352
rect 6167 1302 6220 1318
rect 6250 1488 6306 1512
rect 6250 1454 6261 1488
rect 6295 1454 6306 1488
rect 6250 1420 6306 1454
rect 6250 1386 6261 1420
rect 6295 1386 6306 1420
rect 6250 1352 6306 1386
rect 6250 1318 6261 1352
rect 6295 1318 6306 1352
rect 6250 1302 6306 1318
rect 6336 1488 6389 1512
rect 6336 1454 6347 1488
rect 6381 1454 6389 1488
rect 6336 1420 6389 1454
rect 6336 1386 6347 1420
rect 6381 1386 6389 1420
rect 6336 1352 6389 1386
rect 6336 1318 6347 1352
rect 6381 1318 6389 1352
rect 6336 1302 6389 1318
<< pdiff >>
rect 147 2210 200 2226
rect 147 2176 155 2210
rect 189 2176 200 2210
rect 147 2142 200 2176
rect 147 2108 155 2142
rect 189 2108 200 2142
rect 147 2074 200 2108
rect 147 2040 155 2074
rect 189 2040 200 2074
rect 147 2016 200 2040
rect 230 2210 286 2226
rect 230 2176 241 2210
rect 275 2176 286 2210
rect 230 2142 286 2176
rect 230 2108 241 2142
rect 275 2108 286 2142
rect 230 2074 286 2108
rect 230 2040 241 2074
rect 275 2040 286 2074
rect 230 2016 286 2040
rect 316 2210 372 2226
rect 316 2176 327 2210
rect 361 2176 372 2210
rect 316 2142 372 2176
rect 316 2108 327 2142
rect 361 2108 372 2142
rect 316 2074 372 2108
rect 316 2040 327 2074
rect 361 2040 372 2074
rect 316 2016 372 2040
rect 402 2210 458 2226
rect 402 2176 413 2210
rect 447 2176 458 2210
rect 402 2142 458 2176
rect 402 2108 413 2142
rect 447 2108 458 2142
rect 402 2074 458 2108
rect 402 2040 413 2074
rect 447 2040 458 2074
rect 402 2016 458 2040
rect 488 2210 544 2226
rect 488 2176 499 2210
rect 533 2176 544 2210
rect 488 2142 544 2176
rect 488 2108 499 2142
rect 533 2108 544 2142
rect 488 2074 544 2108
rect 488 2040 499 2074
rect 533 2040 544 2074
rect 488 2016 544 2040
rect 574 2210 630 2226
rect 574 2176 585 2210
rect 619 2176 630 2210
rect 574 2142 630 2176
rect 574 2108 585 2142
rect 619 2108 630 2142
rect 574 2074 630 2108
rect 574 2040 585 2074
rect 619 2040 630 2074
rect 574 2016 630 2040
rect 660 2210 716 2226
rect 660 2176 671 2210
rect 705 2176 716 2210
rect 660 2142 716 2176
rect 660 2108 671 2142
rect 705 2108 716 2142
rect 660 2074 716 2108
rect 660 2040 671 2074
rect 705 2040 716 2074
rect 660 2016 716 2040
rect 746 2210 802 2226
rect 746 2176 757 2210
rect 791 2176 802 2210
rect 746 2142 802 2176
rect 746 2108 757 2142
rect 791 2108 802 2142
rect 746 2074 802 2108
rect 746 2040 757 2074
rect 791 2040 802 2074
rect 746 2016 802 2040
rect 832 2210 888 2226
rect 832 2176 843 2210
rect 877 2176 888 2210
rect 832 2142 888 2176
rect 832 2108 843 2142
rect 877 2108 888 2142
rect 832 2074 888 2108
rect 832 2040 843 2074
rect 877 2040 888 2074
rect 832 2016 888 2040
rect 918 2210 974 2226
rect 918 2176 929 2210
rect 963 2176 974 2210
rect 918 2142 974 2176
rect 918 2108 929 2142
rect 963 2108 974 2142
rect 918 2074 974 2108
rect 918 2040 929 2074
rect 963 2040 974 2074
rect 918 2016 974 2040
rect 1004 2210 1060 2226
rect 1004 2176 1015 2210
rect 1049 2176 1060 2210
rect 1004 2142 1060 2176
rect 1004 2108 1015 2142
rect 1049 2108 1060 2142
rect 1004 2074 1060 2108
rect 1004 2040 1015 2074
rect 1049 2040 1060 2074
rect 1004 2016 1060 2040
rect 1090 2210 1146 2226
rect 1090 2176 1101 2210
rect 1135 2176 1146 2210
rect 1090 2142 1146 2176
rect 1090 2108 1101 2142
rect 1135 2108 1146 2142
rect 1090 2074 1146 2108
rect 1090 2040 1101 2074
rect 1135 2040 1146 2074
rect 1090 2016 1146 2040
rect 1176 2210 1232 2226
rect 1176 2176 1187 2210
rect 1221 2176 1232 2210
rect 1176 2142 1232 2176
rect 1176 2108 1187 2142
rect 1221 2108 1232 2142
rect 1176 2074 1232 2108
rect 1176 2040 1187 2074
rect 1221 2040 1232 2074
rect 1176 2016 1232 2040
rect 1262 2210 1318 2226
rect 1262 2176 1273 2210
rect 1307 2176 1318 2210
rect 1262 2142 1318 2176
rect 1262 2108 1273 2142
rect 1307 2108 1318 2142
rect 1262 2074 1318 2108
rect 1262 2040 1273 2074
rect 1307 2040 1318 2074
rect 1262 2016 1318 2040
rect 1348 2210 1404 2226
rect 1348 2176 1359 2210
rect 1393 2176 1404 2210
rect 1348 2142 1404 2176
rect 1348 2108 1359 2142
rect 1393 2108 1404 2142
rect 1348 2074 1404 2108
rect 1348 2040 1359 2074
rect 1393 2040 1404 2074
rect 1348 2016 1404 2040
rect 1434 2210 1490 2226
rect 1434 2176 1445 2210
rect 1479 2176 1490 2210
rect 1434 2142 1490 2176
rect 1434 2108 1445 2142
rect 1479 2108 1490 2142
rect 1434 2074 1490 2108
rect 1434 2040 1445 2074
rect 1479 2040 1490 2074
rect 1434 2016 1490 2040
rect 1520 2210 1576 2226
rect 1520 2176 1531 2210
rect 1565 2176 1576 2210
rect 1520 2142 1576 2176
rect 1520 2108 1531 2142
rect 1565 2108 1576 2142
rect 1520 2074 1576 2108
rect 1520 2040 1531 2074
rect 1565 2040 1576 2074
rect 1520 2016 1576 2040
rect 1606 2210 1662 2226
rect 1606 2176 1617 2210
rect 1651 2176 1662 2210
rect 1606 2142 1662 2176
rect 1606 2108 1617 2142
rect 1651 2108 1662 2142
rect 1606 2074 1662 2108
rect 1606 2040 1617 2074
rect 1651 2040 1662 2074
rect 1606 2016 1662 2040
rect 1692 2210 1748 2226
rect 1692 2176 1703 2210
rect 1737 2176 1748 2210
rect 1692 2142 1748 2176
rect 1692 2108 1703 2142
rect 1737 2108 1748 2142
rect 1692 2074 1748 2108
rect 1692 2040 1703 2074
rect 1737 2040 1748 2074
rect 1692 2016 1748 2040
rect 1778 2210 1834 2226
rect 1778 2176 1789 2210
rect 1823 2176 1834 2210
rect 1778 2142 1834 2176
rect 1778 2108 1789 2142
rect 1823 2108 1834 2142
rect 1778 2074 1834 2108
rect 1778 2040 1789 2074
rect 1823 2040 1834 2074
rect 1778 2016 1834 2040
rect 1864 2210 1920 2226
rect 1864 2176 1875 2210
rect 1909 2176 1920 2210
rect 1864 2142 1920 2176
rect 1864 2108 1875 2142
rect 1909 2108 1920 2142
rect 1864 2074 1920 2108
rect 1864 2040 1875 2074
rect 1909 2040 1920 2074
rect 1864 2016 1920 2040
rect 1950 2210 2006 2226
rect 1950 2176 1961 2210
rect 1995 2176 2006 2210
rect 1950 2142 2006 2176
rect 1950 2108 1961 2142
rect 1995 2108 2006 2142
rect 1950 2074 2006 2108
rect 1950 2040 1961 2074
rect 1995 2040 2006 2074
rect 1950 2016 2006 2040
rect 2036 2210 2092 2226
rect 2036 2176 2047 2210
rect 2081 2176 2092 2210
rect 2036 2142 2092 2176
rect 2036 2108 2047 2142
rect 2081 2108 2092 2142
rect 2036 2074 2092 2108
rect 2036 2040 2047 2074
rect 2081 2040 2092 2074
rect 2036 2016 2092 2040
rect 2122 2210 2178 2226
rect 2122 2176 2133 2210
rect 2167 2176 2178 2210
rect 2122 2142 2178 2176
rect 2122 2108 2133 2142
rect 2167 2108 2178 2142
rect 2122 2074 2178 2108
rect 2122 2040 2133 2074
rect 2167 2040 2178 2074
rect 2122 2016 2178 2040
rect 2208 2210 2261 2226
rect 2208 2176 2219 2210
rect 2253 2176 2261 2210
rect 2208 2142 2261 2176
rect 2208 2108 2219 2142
rect 2253 2108 2261 2142
rect 2208 2074 2261 2108
rect 2208 2040 2219 2074
rect 2253 2040 2261 2074
rect 2208 2016 2261 2040
rect 2555 2210 2608 2226
rect 2555 2176 2563 2210
rect 2597 2176 2608 2210
rect 2555 2142 2608 2176
rect 2555 2108 2563 2142
rect 2597 2108 2608 2142
rect 2555 2074 2608 2108
rect 2555 2040 2563 2074
rect 2597 2040 2608 2074
rect 2555 2016 2608 2040
rect 2638 2210 2694 2226
rect 2638 2176 2649 2210
rect 2683 2176 2694 2210
rect 2638 2142 2694 2176
rect 2638 2108 2649 2142
rect 2683 2108 2694 2142
rect 2638 2074 2694 2108
rect 2638 2040 2649 2074
rect 2683 2040 2694 2074
rect 2638 2016 2694 2040
rect 2724 2210 2780 2226
rect 2724 2176 2735 2210
rect 2769 2176 2780 2210
rect 2724 2142 2780 2176
rect 2724 2108 2735 2142
rect 2769 2108 2780 2142
rect 2724 2074 2780 2108
rect 2724 2040 2735 2074
rect 2769 2040 2780 2074
rect 2724 2016 2780 2040
rect 2810 2210 2866 2226
rect 2810 2176 2821 2210
rect 2855 2176 2866 2210
rect 2810 2142 2866 2176
rect 2810 2108 2821 2142
rect 2855 2108 2866 2142
rect 2810 2074 2866 2108
rect 2810 2040 2821 2074
rect 2855 2040 2866 2074
rect 2810 2016 2866 2040
rect 2896 2210 2952 2226
rect 2896 2176 2907 2210
rect 2941 2176 2952 2210
rect 2896 2142 2952 2176
rect 2896 2108 2907 2142
rect 2941 2108 2952 2142
rect 2896 2074 2952 2108
rect 2896 2040 2907 2074
rect 2941 2040 2952 2074
rect 2896 2016 2952 2040
rect 2982 2210 3038 2226
rect 2982 2176 2993 2210
rect 3027 2176 3038 2210
rect 2982 2142 3038 2176
rect 2982 2108 2993 2142
rect 3027 2108 3038 2142
rect 2982 2074 3038 2108
rect 2982 2040 2993 2074
rect 3027 2040 3038 2074
rect 2982 2016 3038 2040
rect 3068 2210 3124 2226
rect 3068 2176 3079 2210
rect 3113 2176 3124 2210
rect 3068 2142 3124 2176
rect 3068 2108 3079 2142
rect 3113 2108 3124 2142
rect 3068 2074 3124 2108
rect 3068 2040 3079 2074
rect 3113 2040 3124 2074
rect 3068 2016 3124 2040
rect 3154 2210 3210 2226
rect 3154 2176 3165 2210
rect 3199 2176 3210 2210
rect 3154 2142 3210 2176
rect 3154 2108 3165 2142
rect 3199 2108 3210 2142
rect 3154 2074 3210 2108
rect 3154 2040 3165 2074
rect 3199 2040 3210 2074
rect 3154 2016 3210 2040
rect 3240 2210 3296 2226
rect 3240 2176 3251 2210
rect 3285 2176 3296 2210
rect 3240 2142 3296 2176
rect 3240 2108 3251 2142
rect 3285 2108 3296 2142
rect 3240 2074 3296 2108
rect 3240 2040 3251 2074
rect 3285 2040 3296 2074
rect 3240 2016 3296 2040
rect 3326 2210 3382 2226
rect 3326 2176 3337 2210
rect 3371 2176 3382 2210
rect 3326 2142 3382 2176
rect 3326 2108 3337 2142
rect 3371 2108 3382 2142
rect 3326 2074 3382 2108
rect 3326 2040 3337 2074
rect 3371 2040 3382 2074
rect 3326 2016 3382 2040
rect 3412 2210 3468 2226
rect 3412 2176 3423 2210
rect 3457 2176 3468 2210
rect 3412 2142 3468 2176
rect 3412 2108 3423 2142
rect 3457 2108 3468 2142
rect 3412 2074 3468 2108
rect 3412 2040 3423 2074
rect 3457 2040 3468 2074
rect 3412 2016 3468 2040
rect 3498 2210 3554 2226
rect 3498 2176 3509 2210
rect 3543 2176 3554 2210
rect 3498 2142 3554 2176
rect 3498 2108 3509 2142
rect 3543 2108 3554 2142
rect 3498 2074 3554 2108
rect 3498 2040 3509 2074
rect 3543 2040 3554 2074
rect 3498 2016 3554 2040
rect 3584 2210 3637 2226
rect 3584 2176 3595 2210
rect 3629 2176 3637 2210
rect 3584 2142 3637 2176
rect 3584 2108 3595 2142
rect 3629 2108 3637 2142
rect 3584 2074 3637 2108
rect 3584 2040 3595 2074
rect 3629 2040 3637 2074
rect 6683 2210 6736 2226
rect 6683 2176 6691 2210
rect 6725 2176 6736 2210
rect 6683 2142 6736 2176
rect 6683 2108 6691 2142
rect 6725 2108 6736 2142
rect 6683 2074 6736 2108
rect 3584 2016 3637 2040
rect 6683 2040 6691 2074
rect 6725 2040 6736 2074
rect 6683 2016 6736 2040
rect 6766 2210 6822 2226
rect 6766 2176 6777 2210
rect 6811 2176 6822 2210
rect 6766 2142 6822 2176
rect 6766 2108 6777 2142
rect 6811 2108 6822 2142
rect 6766 2074 6822 2108
rect 6766 2040 6777 2074
rect 6811 2040 6822 2074
rect 6766 2016 6822 2040
rect 6852 2210 6905 2226
rect 6852 2176 6863 2210
rect 6897 2176 6905 2210
rect 6852 2142 6905 2176
rect 6852 2108 6863 2142
rect 6897 2108 6905 2142
rect 6852 2074 6905 2108
rect 6852 2040 6863 2074
rect 6897 2040 6905 2074
rect 6852 2016 6905 2040
rect 7199 2210 7252 2226
rect 7199 2176 7207 2210
rect 7241 2176 7252 2210
rect 7199 2142 7252 2176
rect 7199 2108 7207 2142
rect 7241 2108 7252 2142
rect 7199 2074 7252 2108
rect 7199 2040 7207 2074
rect 7241 2040 7252 2074
rect 7199 2016 7252 2040
rect 7282 2210 7338 2226
rect 7282 2176 7293 2210
rect 7327 2176 7338 2210
rect 7282 2142 7338 2176
rect 7282 2108 7293 2142
rect 7327 2108 7338 2142
rect 7282 2074 7338 2108
rect 7282 2040 7293 2074
rect 7327 2040 7338 2074
rect 7282 2016 7338 2040
rect 7368 2210 7424 2226
rect 7368 2176 7379 2210
rect 7413 2176 7424 2210
rect 7368 2142 7424 2176
rect 7368 2108 7379 2142
rect 7413 2108 7424 2142
rect 7368 2074 7424 2108
rect 7368 2040 7379 2074
rect 7413 2040 7424 2074
rect 7368 2016 7424 2040
rect 7454 2210 7510 2226
rect 7454 2176 7465 2210
rect 7499 2176 7510 2210
rect 7454 2142 7510 2176
rect 7454 2108 7465 2142
rect 7499 2108 7510 2142
rect 7454 2074 7510 2108
rect 7454 2040 7465 2074
rect 7499 2040 7510 2074
rect 7454 2016 7510 2040
rect 7540 2210 7596 2226
rect 7540 2176 7551 2210
rect 7585 2176 7596 2210
rect 7540 2142 7596 2176
rect 7540 2108 7551 2142
rect 7585 2108 7596 2142
rect 7540 2074 7596 2108
rect 7540 2040 7551 2074
rect 7585 2040 7596 2074
rect 7540 2016 7596 2040
rect 7626 2210 7682 2226
rect 7626 2176 7637 2210
rect 7671 2176 7682 2210
rect 7626 2142 7682 2176
rect 7626 2108 7637 2142
rect 7671 2108 7682 2142
rect 7626 2074 7682 2108
rect 7626 2040 7637 2074
rect 7671 2040 7682 2074
rect 7626 2016 7682 2040
rect 7712 2210 7768 2226
rect 7712 2176 7723 2210
rect 7757 2176 7768 2210
rect 7712 2142 7768 2176
rect 7712 2108 7723 2142
rect 7757 2108 7768 2142
rect 7712 2074 7768 2108
rect 7712 2040 7723 2074
rect 7757 2040 7768 2074
rect 7712 2016 7768 2040
rect 7798 2210 7854 2226
rect 7798 2176 7809 2210
rect 7843 2176 7854 2210
rect 7798 2142 7854 2176
rect 7798 2108 7809 2142
rect 7843 2108 7854 2142
rect 7798 2074 7854 2108
rect 7798 2040 7809 2074
rect 7843 2040 7854 2074
rect 7798 2016 7854 2040
rect 7884 2210 7940 2226
rect 7884 2176 7895 2210
rect 7929 2176 7940 2210
rect 7884 2142 7940 2176
rect 7884 2108 7895 2142
rect 7929 2108 7940 2142
rect 7884 2074 7940 2108
rect 7884 2040 7895 2074
rect 7929 2040 7940 2074
rect 7884 2016 7940 2040
rect 7970 2210 8026 2226
rect 7970 2176 7981 2210
rect 8015 2176 8026 2210
rect 7970 2142 8026 2176
rect 7970 2108 7981 2142
rect 8015 2108 8026 2142
rect 7970 2074 8026 2108
rect 7970 2040 7981 2074
rect 8015 2040 8026 2074
rect 7970 2016 8026 2040
rect 8056 2210 8112 2226
rect 8056 2176 8067 2210
rect 8101 2176 8112 2210
rect 8056 2142 8112 2176
rect 8056 2108 8067 2142
rect 8101 2108 8112 2142
rect 8056 2074 8112 2108
rect 8056 2040 8067 2074
rect 8101 2040 8112 2074
rect 8056 2016 8112 2040
rect 8142 2210 8198 2226
rect 8142 2176 8153 2210
rect 8187 2176 8198 2210
rect 8142 2142 8198 2176
rect 8142 2108 8153 2142
rect 8187 2108 8198 2142
rect 8142 2074 8198 2108
rect 8142 2040 8153 2074
rect 8187 2040 8198 2074
rect 8142 2016 8198 2040
rect 8228 2210 8284 2226
rect 8228 2176 8239 2210
rect 8273 2176 8284 2210
rect 8228 2142 8284 2176
rect 8228 2108 8239 2142
rect 8273 2108 8284 2142
rect 8228 2074 8284 2108
rect 8228 2040 8239 2074
rect 8273 2040 8284 2074
rect 8228 2016 8284 2040
rect 8314 2210 8370 2226
rect 8314 2176 8325 2210
rect 8359 2176 8370 2210
rect 8314 2142 8370 2176
rect 8314 2108 8325 2142
rect 8359 2108 8370 2142
rect 8314 2074 8370 2108
rect 8314 2040 8325 2074
rect 8359 2040 8370 2074
rect 8314 2016 8370 2040
rect 8400 2210 8456 2226
rect 8400 2176 8411 2210
rect 8445 2176 8456 2210
rect 8400 2142 8456 2176
rect 8400 2108 8411 2142
rect 8445 2108 8456 2142
rect 8400 2074 8456 2108
rect 8400 2040 8411 2074
rect 8445 2040 8456 2074
rect 8400 2016 8456 2040
rect 8486 2210 8542 2226
rect 8486 2176 8497 2210
rect 8531 2176 8542 2210
rect 8486 2142 8542 2176
rect 8486 2108 8497 2142
rect 8531 2108 8542 2142
rect 8486 2074 8542 2108
rect 8486 2040 8497 2074
rect 8531 2040 8542 2074
rect 8486 2016 8542 2040
rect 8572 2210 8628 2226
rect 8572 2176 8583 2210
rect 8617 2176 8628 2210
rect 8572 2142 8628 2176
rect 8572 2108 8583 2142
rect 8617 2108 8628 2142
rect 8572 2074 8628 2108
rect 8572 2040 8583 2074
rect 8617 2040 8628 2074
rect 8572 2016 8628 2040
rect 8658 2210 8714 2226
rect 8658 2176 8669 2210
rect 8703 2176 8714 2210
rect 8658 2142 8714 2176
rect 8658 2108 8669 2142
rect 8703 2108 8714 2142
rect 8658 2074 8714 2108
rect 8658 2040 8669 2074
rect 8703 2040 8714 2074
rect 8658 2016 8714 2040
rect 8744 2210 8800 2226
rect 8744 2176 8755 2210
rect 8789 2176 8800 2210
rect 8744 2142 8800 2176
rect 8744 2108 8755 2142
rect 8789 2108 8800 2142
rect 8744 2074 8800 2108
rect 8744 2040 8755 2074
rect 8789 2040 8800 2074
rect 8744 2016 8800 2040
rect 8830 2210 8886 2226
rect 8830 2176 8841 2210
rect 8875 2176 8886 2210
rect 8830 2142 8886 2176
rect 8830 2108 8841 2142
rect 8875 2108 8886 2142
rect 8830 2074 8886 2108
rect 8830 2040 8841 2074
rect 8875 2040 8886 2074
rect 8830 2016 8886 2040
rect 8916 2210 8972 2226
rect 8916 2176 8927 2210
rect 8961 2176 8972 2210
rect 8916 2142 8972 2176
rect 8916 2108 8927 2142
rect 8961 2108 8972 2142
rect 8916 2074 8972 2108
rect 8916 2040 8927 2074
rect 8961 2040 8972 2074
rect 8916 2016 8972 2040
rect 9002 2210 9058 2226
rect 9002 2176 9013 2210
rect 9047 2176 9058 2210
rect 9002 2142 9058 2176
rect 9002 2108 9013 2142
rect 9047 2108 9058 2142
rect 9002 2074 9058 2108
rect 9002 2040 9013 2074
rect 9047 2040 9058 2074
rect 9002 2016 9058 2040
rect 9088 2210 9144 2226
rect 9088 2176 9099 2210
rect 9133 2176 9144 2210
rect 9088 2142 9144 2176
rect 9088 2108 9099 2142
rect 9133 2108 9144 2142
rect 9088 2074 9144 2108
rect 9088 2040 9099 2074
rect 9133 2040 9144 2074
rect 9088 2016 9144 2040
rect 9174 2210 9230 2226
rect 9174 2176 9185 2210
rect 9219 2176 9230 2210
rect 9174 2142 9230 2176
rect 9174 2108 9185 2142
rect 9219 2108 9230 2142
rect 9174 2074 9230 2108
rect 9174 2040 9185 2074
rect 9219 2040 9230 2074
rect 9174 2016 9230 2040
rect 9260 2210 9316 2226
rect 9260 2176 9271 2210
rect 9305 2176 9316 2210
rect 9260 2142 9316 2176
rect 9260 2108 9271 2142
rect 9305 2108 9316 2142
rect 9260 2074 9316 2108
rect 9260 2040 9271 2074
rect 9305 2040 9316 2074
rect 9260 2016 9316 2040
rect 9346 2210 9402 2226
rect 9346 2176 9357 2210
rect 9391 2176 9402 2210
rect 9346 2142 9402 2176
rect 9346 2108 9357 2142
rect 9391 2108 9402 2142
rect 9346 2074 9402 2108
rect 9346 2040 9357 2074
rect 9391 2040 9402 2074
rect 9346 2016 9402 2040
rect 9432 2210 9488 2226
rect 9432 2176 9443 2210
rect 9477 2176 9488 2210
rect 9432 2142 9488 2176
rect 9432 2108 9443 2142
rect 9477 2108 9488 2142
rect 9432 2074 9488 2108
rect 9432 2040 9443 2074
rect 9477 2040 9488 2074
rect 9432 2016 9488 2040
rect 9518 2210 9574 2226
rect 9518 2176 9529 2210
rect 9563 2176 9574 2210
rect 9518 2142 9574 2176
rect 9518 2108 9529 2142
rect 9563 2108 9574 2142
rect 9518 2074 9574 2108
rect 9518 2040 9529 2074
rect 9563 2040 9574 2074
rect 9518 2016 9574 2040
rect 9604 2210 9660 2226
rect 9604 2176 9615 2210
rect 9649 2176 9660 2210
rect 9604 2142 9660 2176
rect 9604 2108 9615 2142
rect 9649 2108 9660 2142
rect 9604 2074 9660 2108
rect 9604 2040 9615 2074
rect 9649 2040 9660 2074
rect 9604 2016 9660 2040
rect 9690 2210 9746 2226
rect 9690 2176 9701 2210
rect 9735 2176 9746 2210
rect 9690 2142 9746 2176
rect 9690 2108 9701 2142
rect 9735 2108 9746 2142
rect 9690 2074 9746 2108
rect 9690 2040 9701 2074
rect 9735 2040 9746 2074
rect 9690 2016 9746 2040
rect 9776 2210 9832 2226
rect 9776 2176 9787 2210
rect 9821 2176 9832 2210
rect 9776 2142 9832 2176
rect 9776 2108 9787 2142
rect 9821 2108 9832 2142
rect 9776 2074 9832 2108
rect 9776 2040 9787 2074
rect 9821 2040 9832 2074
rect 9776 2016 9832 2040
rect 9862 2210 9918 2226
rect 9862 2176 9873 2210
rect 9907 2176 9918 2210
rect 9862 2142 9918 2176
rect 9862 2108 9873 2142
rect 9907 2108 9918 2142
rect 9862 2074 9918 2108
rect 9862 2040 9873 2074
rect 9907 2040 9918 2074
rect 9862 2016 9918 2040
rect 9948 2210 10004 2226
rect 9948 2176 9959 2210
rect 9993 2176 10004 2210
rect 9948 2142 10004 2176
rect 9948 2108 9959 2142
rect 9993 2108 10004 2142
rect 9948 2074 10004 2108
rect 9948 2040 9959 2074
rect 9993 2040 10004 2074
rect 9948 2016 10004 2040
rect 10034 2210 10090 2226
rect 10034 2176 10045 2210
rect 10079 2176 10090 2210
rect 10034 2142 10090 2176
rect 10034 2108 10045 2142
rect 10079 2108 10090 2142
rect 10034 2074 10090 2108
rect 10034 2040 10045 2074
rect 10079 2040 10090 2074
rect 10034 2016 10090 2040
rect 10120 2210 10176 2226
rect 10120 2176 10131 2210
rect 10165 2176 10176 2210
rect 10120 2142 10176 2176
rect 10120 2108 10131 2142
rect 10165 2108 10176 2142
rect 10120 2074 10176 2108
rect 10120 2040 10131 2074
rect 10165 2040 10176 2074
rect 10120 2016 10176 2040
rect 10206 2210 10262 2226
rect 10206 2176 10217 2210
rect 10251 2176 10262 2210
rect 10206 2142 10262 2176
rect 10206 2108 10217 2142
rect 10251 2108 10262 2142
rect 10206 2074 10262 2108
rect 10206 2040 10217 2074
rect 10251 2040 10262 2074
rect 10206 2016 10262 2040
rect 10292 2210 10348 2226
rect 10292 2176 10303 2210
rect 10337 2176 10348 2210
rect 10292 2142 10348 2176
rect 10292 2108 10303 2142
rect 10337 2108 10348 2142
rect 10292 2074 10348 2108
rect 10292 2040 10303 2074
rect 10337 2040 10348 2074
rect 10292 2016 10348 2040
rect 10378 2210 10434 2226
rect 10378 2176 10389 2210
rect 10423 2176 10434 2210
rect 10378 2142 10434 2176
rect 10378 2108 10389 2142
rect 10423 2108 10434 2142
rect 10378 2074 10434 2108
rect 10378 2040 10389 2074
rect 10423 2040 10434 2074
rect 10378 2016 10434 2040
rect 10464 2210 10520 2226
rect 10464 2176 10475 2210
rect 10509 2176 10520 2210
rect 10464 2142 10520 2176
rect 10464 2108 10475 2142
rect 10509 2108 10520 2142
rect 10464 2074 10520 2108
rect 10464 2040 10475 2074
rect 10509 2040 10520 2074
rect 10464 2016 10520 2040
rect 10550 2210 10606 2226
rect 10550 2176 10561 2210
rect 10595 2176 10606 2210
rect 10550 2142 10606 2176
rect 10550 2108 10561 2142
rect 10595 2108 10606 2142
rect 10550 2074 10606 2108
rect 10550 2040 10561 2074
rect 10595 2040 10606 2074
rect 10550 2016 10606 2040
rect 10636 2210 10692 2226
rect 10636 2176 10647 2210
rect 10681 2176 10692 2210
rect 10636 2142 10692 2176
rect 10636 2108 10647 2142
rect 10681 2108 10692 2142
rect 10636 2074 10692 2108
rect 10636 2040 10647 2074
rect 10681 2040 10692 2074
rect 10636 2016 10692 2040
rect 10722 2210 10778 2226
rect 10722 2176 10733 2210
rect 10767 2176 10778 2210
rect 10722 2142 10778 2176
rect 10722 2108 10733 2142
rect 10767 2108 10778 2142
rect 10722 2074 10778 2108
rect 10722 2040 10733 2074
rect 10767 2040 10778 2074
rect 10722 2016 10778 2040
rect 10808 2210 10864 2226
rect 10808 2176 10819 2210
rect 10853 2176 10864 2210
rect 10808 2142 10864 2176
rect 10808 2108 10819 2142
rect 10853 2108 10864 2142
rect 10808 2074 10864 2108
rect 10808 2040 10819 2074
rect 10853 2040 10864 2074
rect 10808 2016 10864 2040
rect 10894 2210 10950 2226
rect 10894 2176 10905 2210
rect 10939 2176 10950 2210
rect 10894 2142 10950 2176
rect 10894 2108 10905 2142
rect 10939 2108 10950 2142
rect 10894 2074 10950 2108
rect 10894 2040 10905 2074
rect 10939 2040 10950 2074
rect 10894 2016 10950 2040
rect 10980 2210 11036 2226
rect 10980 2176 10991 2210
rect 11025 2176 11036 2210
rect 10980 2142 11036 2176
rect 10980 2108 10991 2142
rect 11025 2108 11036 2142
rect 10980 2074 11036 2108
rect 10980 2040 10991 2074
rect 11025 2040 11036 2074
rect 10980 2016 11036 2040
rect 11066 2210 11122 2226
rect 11066 2176 11077 2210
rect 11111 2176 11122 2210
rect 11066 2142 11122 2176
rect 11066 2108 11077 2142
rect 11111 2108 11122 2142
rect 11066 2074 11122 2108
rect 11066 2040 11077 2074
rect 11111 2040 11122 2074
rect 11066 2016 11122 2040
rect 11152 2210 11208 2226
rect 11152 2176 11163 2210
rect 11197 2176 11208 2210
rect 11152 2142 11208 2176
rect 11152 2108 11163 2142
rect 11197 2108 11208 2142
rect 11152 2074 11208 2108
rect 11152 2040 11163 2074
rect 11197 2040 11208 2074
rect 11152 2016 11208 2040
rect 11238 2210 11294 2226
rect 11238 2176 11249 2210
rect 11283 2176 11294 2210
rect 11238 2142 11294 2176
rect 11238 2108 11249 2142
rect 11283 2108 11294 2142
rect 11238 2074 11294 2108
rect 11238 2040 11249 2074
rect 11283 2040 11294 2074
rect 11238 2016 11294 2040
rect 11324 2210 11377 2226
rect 11324 2176 11335 2210
rect 11369 2176 11377 2210
rect 11324 2142 11377 2176
rect 11324 2108 11335 2142
rect 11369 2108 11377 2142
rect 11324 2074 11377 2108
rect 11324 2040 11335 2074
rect 11369 2040 11377 2074
rect 11324 2016 11377 2040
rect 3931 1454 3984 1470
rect 3931 1420 3939 1454
rect 3973 1420 3984 1454
rect 3931 1386 3984 1420
rect 3931 1352 3939 1386
rect 3973 1352 3984 1386
rect 3931 1318 3984 1352
rect 3931 1284 3939 1318
rect 3973 1284 3984 1318
rect 3931 1260 3984 1284
rect 4014 1454 4070 1470
rect 4014 1420 4025 1454
rect 4059 1420 4070 1454
rect 4014 1386 4070 1420
rect 4014 1352 4025 1386
rect 4059 1352 4070 1386
rect 4014 1318 4070 1352
rect 4014 1284 4025 1318
rect 4059 1284 4070 1318
rect 4014 1260 4070 1284
rect 4100 1454 4156 1470
rect 4100 1420 4111 1454
rect 4145 1420 4156 1454
rect 4100 1386 4156 1420
rect 4100 1352 4111 1386
rect 4145 1352 4156 1386
rect 4100 1318 4156 1352
rect 4100 1284 4111 1318
rect 4145 1284 4156 1318
rect 4100 1260 4156 1284
rect 4186 1454 4242 1470
rect 4186 1420 4197 1454
rect 4231 1420 4242 1454
rect 4186 1386 4242 1420
rect 4186 1352 4197 1386
rect 4231 1352 4242 1386
rect 4186 1318 4242 1352
rect 4186 1284 4197 1318
rect 4231 1284 4242 1318
rect 4186 1260 4242 1284
rect 4272 1454 4328 1470
rect 4272 1420 4283 1454
rect 4317 1420 4328 1454
rect 4272 1386 4328 1420
rect 4272 1352 4283 1386
rect 4317 1352 4328 1386
rect 4272 1318 4328 1352
rect 4272 1284 4283 1318
rect 4317 1284 4328 1318
rect 4272 1260 4328 1284
rect 4358 1454 4414 1470
rect 4358 1420 4369 1454
rect 4403 1420 4414 1454
rect 4358 1386 4414 1420
rect 4358 1352 4369 1386
rect 4403 1352 4414 1386
rect 4358 1318 4414 1352
rect 4358 1284 4369 1318
rect 4403 1284 4414 1318
rect 4358 1260 4414 1284
rect 4444 1454 4500 1470
rect 4444 1420 4455 1454
rect 4489 1420 4500 1454
rect 4444 1386 4500 1420
rect 4444 1352 4455 1386
rect 4489 1352 4500 1386
rect 4444 1318 4500 1352
rect 4444 1284 4455 1318
rect 4489 1284 4500 1318
rect 4444 1260 4500 1284
rect 4530 1454 4586 1470
rect 4530 1420 4541 1454
rect 4575 1420 4586 1454
rect 4530 1386 4586 1420
rect 4530 1352 4541 1386
rect 4575 1352 4586 1386
rect 4530 1318 4586 1352
rect 4530 1284 4541 1318
rect 4575 1284 4586 1318
rect 4530 1260 4586 1284
rect 4616 1454 4672 1470
rect 4616 1420 4627 1454
rect 4661 1420 4672 1454
rect 4616 1386 4672 1420
rect 4616 1352 4627 1386
rect 4661 1352 4672 1386
rect 4616 1318 4672 1352
rect 4616 1284 4627 1318
rect 4661 1284 4672 1318
rect 4616 1260 4672 1284
rect 4702 1454 4758 1470
rect 4702 1420 4713 1454
rect 4747 1420 4758 1454
rect 4702 1386 4758 1420
rect 4702 1352 4713 1386
rect 4747 1352 4758 1386
rect 4702 1318 4758 1352
rect 4702 1284 4713 1318
rect 4747 1284 4758 1318
rect 4702 1260 4758 1284
rect 4788 1454 4844 1470
rect 4788 1420 4799 1454
rect 4833 1420 4844 1454
rect 4788 1386 4844 1420
rect 4788 1352 4799 1386
rect 4833 1352 4844 1386
rect 4788 1318 4844 1352
rect 4788 1284 4799 1318
rect 4833 1284 4844 1318
rect 4788 1260 4844 1284
rect 4874 1454 4930 1470
rect 4874 1420 4885 1454
rect 4919 1420 4930 1454
rect 4874 1386 4930 1420
rect 4874 1352 4885 1386
rect 4919 1352 4930 1386
rect 4874 1318 4930 1352
rect 4874 1284 4885 1318
rect 4919 1284 4930 1318
rect 4874 1260 4930 1284
rect 4960 1454 5013 1470
rect 4960 1420 4971 1454
rect 5005 1420 5013 1454
rect 4960 1386 5013 1420
rect 4960 1352 4971 1386
rect 5005 1352 5013 1386
rect 4960 1318 5013 1352
rect 4960 1284 4971 1318
rect 5005 1284 5013 1318
rect 4960 1260 5013 1284
rect 5307 1454 5360 1470
rect 5307 1420 5315 1454
rect 5349 1420 5360 1454
rect 5307 1386 5360 1420
rect 5307 1352 5315 1386
rect 5349 1352 5360 1386
rect 5307 1318 5360 1352
rect 5307 1284 5315 1318
rect 5349 1284 5360 1318
rect 5307 1260 5360 1284
rect 5390 1454 5446 1470
rect 5390 1420 5401 1454
rect 5435 1420 5446 1454
rect 5390 1386 5446 1420
rect 5390 1352 5401 1386
rect 5435 1352 5446 1386
rect 5390 1318 5446 1352
rect 5390 1284 5401 1318
rect 5435 1284 5446 1318
rect 5390 1260 5446 1284
rect 5476 1454 5532 1470
rect 5476 1420 5487 1454
rect 5521 1420 5532 1454
rect 5476 1386 5532 1420
rect 5476 1352 5487 1386
rect 5521 1352 5532 1386
rect 5476 1318 5532 1352
rect 5476 1284 5487 1318
rect 5521 1284 5532 1318
rect 5476 1260 5532 1284
rect 5562 1454 5618 1470
rect 5562 1420 5573 1454
rect 5607 1420 5618 1454
rect 5562 1386 5618 1420
rect 5562 1352 5573 1386
rect 5607 1352 5618 1386
rect 5562 1318 5618 1352
rect 5562 1284 5573 1318
rect 5607 1284 5618 1318
rect 5562 1260 5618 1284
rect 5648 1454 5704 1470
rect 5648 1420 5659 1454
rect 5693 1420 5704 1454
rect 5648 1386 5704 1420
rect 5648 1352 5659 1386
rect 5693 1352 5704 1386
rect 5648 1318 5704 1352
rect 5648 1284 5659 1318
rect 5693 1284 5704 1318
rect 5648 1260 5704 1284
rect 5734 1454 5790 1470
rect 5734 1420 5745 1454
rect 5779 1420 5790 1454
rect 5734 1386 5790 1420
rect 5734 1352 5745 1386
rect 5779 1352 5790 1386
rect 5734 1318 5790 1352
rect 5734 1284 5745 1318
rect 5779 1284 5790 1318
rect 5734 1260 5790 1284
rect 5820 1454 5873 1470
rect 5820 1420 5831 1454
rect 5865 1420 5873 1454
rect 5820 1386 5873 1420
rect 5820 1352 5831 1386
rect 5865 1352 5873 1386
rect 5820 1318 5873 1352
rect 5820 1284 5831 1318
rect 5865 1284 5873 1318
rect 5820 1260 5873 1284
rect 147 1034 200 1050
rect 147 1000 155 1034
rect 189 1000 200 1034
rect 147 966 200 1000
rect 147 932 155 966
rect 189 932 200 966
rect 147 898 200 932
rect 147 864 155 898
rect 189 864 200 898
rect 147 840 200 864
rect 230 1034 286 1050
rect 230 1000 241 1034
rect 275 1000 286 1034
rect 230 966 286 1000
rect 230 932 241 966
rect 275 932 286 966
rect 230 898 286 932
rect 230 864 241 898
rect 275 864 286 898
rect 230 840 286 864
rect 316 1034 372 1050
rect 316 1000 327 1034
rect 361 1000 372 1034
rect 316 966 372 1000
rect 316 932 327 966
rect 361 932 372 966
rect 316 898 372 932
rect 316 864 327 898
rect 361 864 372 898
rect 316 840 372 864
rect 402 1034 458 1050
rect 402 1000 413 1034
rect 447 1000 458 1034
rect 402 966 458 1000
rect 402 932 413 966
rect 447 932 458 966
rect 402 898 458 932
rect 402 864 413 898
rect 447 864 458 898
rect 402 840 458 864
rect 488 1034 544 1050
rect 488 1000 499 1034
rect 533 1000 544 1034
rect 488 966 544 1000
rect 488 932 499 966
rect 533 932 544 966
rect 488 898 544 932
rect 488 864 499 898
rect 533 864 544 898
rect 488 840 544 864
rect 574 1034 630 1050
rect 574 1000 585 1034
rect 619 1000 630 1034
rect 574 966 630 1000
rect 574 932 585 966
rect 619 932 630 966
rect 574 898 630 932
rect 574 864 585 898
rect 619 864 630 898
rect 574 840 630 864
rect 660 1034 716 1050
rect 660 1000 671 1034
rect 705 1000 716 1034
rect 660 966 716 1000
rect 660 932 671 966
rect 705 932 716 966
rect 660 898 716 932
rect 660 864 671 898
rect 705 864 716 898
rect 660 840 716 864
rect 746 1034 802 1050
rect 746 1000 757 1034
rect 791 1000 802 1034
rect 746 966 802 1000
rect 746 932 757 966
rect 791 932 802 966
rect 746 898 802 932
rect 746 864 757 898
rect 791 864 802 898
rect 746 840 802 864
rect 832 1034 888 1050
rect 832 1000 843 1034
rect 877 1000 888 1034
rect 832 966 888 1000
rect 832 932 843 966
rect 877 932 888 966
rect 832 898 888 932
rect 832 864 843 898
rect 877 864 888 898
rect 832 840 888 864
rect 918 1034 974 1050
rect 918 1000 929 1034
rect 963 1000 974 1034
rect 918 966 974 1000
rect 918 932 929 966
rect 963 932 974 966
rect 918 898 974 932
rect 918 864 929 898
rect 963 864 974 898
rect 918 840 974 864
rect 1004 1034 1060 1050
rect 1004 1000 1015 1034
rect 1049 1000 1060 1034
rect 1004 966 1060 1000
rect 1004 932 1015 966
rect 1049 932 1060 966
rect 1004 898 1060 932
rect 1004 864 1015 898
rect 1049 864 1060 898
rect 1004 840 1060 864
rect 1090 1034 1146 1050
rect 1090 1000 1101 1034
rect 1135 1000 1146 1034
rect 1090 966 1146 1000
rect 1090 932 1101 966
rect 1135 932 1146 966
rect 1090 898 1146 932
rect 1090 864 1101 898
rect 1135 864 1146 898
rect 1090 840 1146 864
rect 1176 1034 1232 1050
rect 1176 1000 1187 1034
rect 1221 1000 1232 1034
rect 1176 966 1232 1000
rect 1176 932 1187 966
rect 1221 932 1232 966
rect 1176 898 1232 932
rect 1176 864 1187 898
rect 1221 864 1232 898
rect 1176 840 1232 864
rect 1262 1034 1318 1050
rect 1262 1000 1273 1034
rect 1307 1000 1318 1034
rect 1262 966 1318 1000
rect 1262 932 1273 966
rect 1307 932 1318 966
rect 1262 898 1318 932
rect 1262 864 1273 898
rect 1307 864 1318 898
rect 1262 840 1318 864
rect 1348 1034 1404 1050
rect 1348 1000 1359 1034
rect 1393 1000 1404 1034
rect 1348 966 1404 1000
rect 1348 932 1359 966
rect 1393 932 1404 966
rect 1348 898 1404 932
rect 1348 864 1359 898
rect 1393 864 1404 898
rect 1348 840 1404 864
rect 1434 1034 1490 1050
rect 1434 1000 1445 1034
rect 1479 1000 1490 1034
rect 1434 966 1490 1000
rect 1434 932 1445 966
rect 1479 932 1490 966
rect 1434 898 1490 932
rect 1434 864 1445 898
rect 1479 864 1490 898
rect 1434 840 1490 864
rect 1520 1034 1576 1050
rect 1520 1000 1531 1034
rect 1565 1000 1576 1034
rect 1520 966 1576 1000
rect 1520 932 1531 966
rect 1565 932 1576 966
rect 1520 898 1576 932
rect 1520 864 1531 898
rect 1565 864 1576 898
rect 1520 840 1576 864
rect 1606 1034 1662 1050
rect 1606 1000 1617 1034
rect 1651 1000 1662 1034
rect 1606 966 1662 1000
rect 1606 932 1617 966
rect 1651 932 1662 966
rect 1606 898 1662 932
rect 1606 864 1617 898
rect 1651 864 1662 898
rect 1606 840 1662 864
rect 1692 1034 1748 1050
rect 1692 1000 1703 1034
rect 1737 1000 1748 1034
rect 1692 966 1748 1000
rect 1692 932 1703 966
rect 1737 932 1748 966
rect 1692 898 1748 932
rect 1692 864 1703 898
rect 1737 864 1748 898
rect 1692 840 1748 864
rect 1778 1034 1834 1050
rect 1778 1000 1789 1034
rect 1823 1000 1834 1034
rect 1778 966 1834 1000
rect 1778 932 1789 966
rect 1823 932 1834 966
rect 1778 898 1834 932
rect 1778 864 1789 898
rect 1823 864 1834 898
rect 1778 840 1834 864
rect 1864 1034 1920 1050
rect 1864 1000 1875 1034
rect 1909 1000 1920 1034
rect 1864 966 1920 1000
rect 1864 932 1875 966
rect 1909 932 1920 966
rect 1864 898 1920 932
rect 1864 864 1875 898
rect 1909 864 1920 898
rect 1864 840 1920 864
rect 1950 1034 2006 1050
rect 1950 1000 1961 1034
rect 1995 1000 2006 1034
rect 1950 966 2006 1000
rect 1950 932 1961 966
rect 1995 932 2006 966
rect 1950 898 2006 932
rect 1950 864 1961 898
rect 1995 864 2006 898
rect 1950 840 2006 864
rect 2036 1034 2092 1050
rect 2036 1000 2047 1034
rect 2081 1000 2092 1034
rect 2036 966 2092 1000
rect 2036 932 2047 966
rect 2081 932 2092 966
rect 2036 898 2092 932
rect 2036 864 2047 898
rect 2081 864 2092 898
rect 2036 840 2092 864
rect 2122 1034 2178 1050
rect 2122 1000 2133 1034
rect 2167 1000 2178 1034
rect 2122 966 2178 1000
rect 2122 932 2133 966
rect 2167 932 2178 966
rect 2122 898 2178 932
rect 2122 864 2133 898
rect 2167 864 2178 898
rect 2122 840 2178 864
rect 2208 1034 2261 1050
rect 2208 1000 2219 1034
rect 2253 1000 2261 1034
rect 2208 966 2261 1000
rect 2208 932 2219 966
rect 2253 932 2261 966
rect 2208 898 2261 932
rect 2208 864 2219 898
rect 2253 864 2261 898
rect 2208 840 2261 864
rect 2555 1034 2608 1050
rect 2555 1000 2563 1034
rect 2597 1000 2608 1034
rect 2555 966 2608 1000
rect 2555 932 2563 966
rect 2597 932 2608 966
rect 2555 898 2608 932
rect 2555 864 2563 898
rect 2597 864 2608 898
rect 2555 840 2608 864
rect 2638 1034 2694 1050
rect 2638 1000 2649 1034
rect 2683 1000 2694 1034
rect 2638 966 2694 1000
rect 2638 932 2649 966
rect 2683 932 2694 966
rect 2638 898 2694 932
rect 2638 864 2649 898
rect 2683 864 2694 898
rect 2638 840 2694 864
rect 2724 1034 2780 1050
rect 2724 1000 2735 1034
rect 2769 1000 2780 1034
rect 2724 966 2780 1000
rect 2724 932 2735 966
rect 2769 932 2780 966
rect 2724 898 2780 932
rect 2724 864 2735 898
rect 2769 864 2780 898
rect 2724 840 2780 864
rect 2810 1034 2866 1050
rect 2810 1000 2821 1034
rect 2855 1000 2866 1034
rect 2810 966 2866 1000
rect 2810 932 2821 966
rect 2855 932 2866 966
rect 2810 898 2866 932
rect 2810 864 2821 898
rect 2855 864 2866 898
rect 2810 840 2866 864
rect 2896 1034 2952 1050
rect 2896 1000 2907 1034
rect 2941 1000 2952 1034
rect 2896 966 2952 1000
rect 2896 932 2907 966
rect 2941 932 2952 966
rect 2896 898 2952 932
rect 2896 864 2907 898
rect 2941 864 2952 898
rect 2896 840 2952 864
rect 2982 1034 3038 1050
rect 2982 1000 2993 1034
rect 3027 1000 3038 1034
rect 2982 966 3038 1000
rect 2982 932 2993 966
rect 3027 932 3038 966
rect 2982 898 3038 932
rect 2982 864 2993 898
rect 3027 864 3038 898
rect 2982 840 3038 864
rect 3068 1034 3124 1050
rect 3068 1000 3079 1034
rect 3113 1000 3124 1034
rect 3068 966 3124 1000
rect 3068 932 3079 966
rect 3113 932 3124 966
rect 3068 898 3124 932
rect 3068 864 3079 898
rect 3113 864 3124 898
rect 3068 840 3124 864
rect 3154 1034 3210 1050
rect 3154 1000 3165 1034
rect 3199 1000 3210 1034
rect 3154 966 3210 1000
rect 3154 932 3165 966
rect 3199 932 3210 966
rect 3154 898 3210 932
rect 3154 864 3165 898
rect 3199 864 3210 898
rect 3154 840 3210 864
rect 3240 1034 3296 1050
rect 3240 1000 3251 1034
rect 3285 1000 3296 1034
rect 3240 966 3296 1000
rect 3240 932 3251 966
rect 3285 932 3296 966
rect 3240 898 3296 932
rect 3240 864 3251 898
rect 3285 864 3296 898
rect 3240 840 3296 864
rect 3326 1034 3382 1050
rect 3326 1000 3337 1034
rect 3371 1000 3382 1034
rect 3326 966 3382 1000
rect 3326 932 3337 966
rect 3371 932 3382 966
rect 3326 898 3382 932
rect 3326 864 3337 898
rect 3371 864 3382 898
rect 3326 840 3382 864
rect 3412 1034 3468 1050
rect 3412 1000 3423 1034
rect 3457 1000 3468 1034
rect 3412 966 3468 1000
rect 3412 932 3423 966
rect 3457 932 3468 966
rect 3412 898 3468 932
rect 3412 864 3423 898
rect 3457 864 3468 898
rect 3412 840 3468 864
rect 3498 1034 3554 1050
rect 3498 1000 3509 1034
rect 3543 1000 3554 1034
rect 3498 966 3554 1000
rect 3498 932 3509 966
rect 3543 932 3554 966
rect 3498 898 3554 932
rect 3498 864 3509 898
rect 3543 864 3554 898
rect 3498 840 3554 864
rect 3584 1034 3637 1050
rect 3584 1000 3595 1034
rect 3629 1000 3637 1034
rect 3584 966 3637 1000
rect 7199 1034 7252 1050
rect 7199 1000 7207 1034
rect 7241 1000 7252 1034
rect 3584 932 3595 966
rect 3629 932 3637 966
rect 3584 898 3637 932
rect 3584 864 3595 898
rect 3629 864 3637 898
rect 3584 840 3637 864
rect 7199 966 7252 1000
rect 7199 932 7207 966
rect 7241 932 7252 966
rect 7199 898 7252 932
rect 7199 864 7207 898
rect 7241 864 7252 898
rect 7199 840 7252 864
rect 7282 1034 7338 1050
rect 7282 1000 7293 1034
rect 7327 1000 7338 1034
rect 7282 966 7338 1000
rect 7282 932 7293 966
rect 7327 932 7338 966
rect 7282 898 7338 932
rect 7282 864 7293 898
rect 7327 864 7338 898
rect 7282 840 7338 864
rect 7368 1034 7424 1050
rect 7368 1000 7379 1034
rect 7413 1000 7424 1034
rect 7368 966 7424 1000
rect 7368 932 7379 966
rect 7413 932 7424 966
rect 7368 898 7424 932
rect 7368 864 7379 898
rect 7413 864 7424 898
rect 7368 840 7424 864
rect 7454 1034 7510 1050
rect 7454 1000 7465 1034
rect 7499 1000 7510 1034
rect 7454 966 7510 1000
rect 7454 932 7465 966
rect 7499 932 7510 966
rect 7454 898 7510 932
rect 7454 864 7465 898
rect 7499 864 7510 898
rect 7454 840 7510 864
rect 7540 1034 7596 1050
rect 7540 1000 7551 1034
rect 7585 1000 7596 1034
rect 7540 966 7596 1000
rect 7540 932 7551 966
rect 7585 932 7596 966
rect 7540 898 7596 932
rect 7540 864 7551 898
rect 7585 864 7596 898
rect 7540 840 7596 864
rect 7626 1034 7682 1050
rect 7626 1000 7637 1034
rect 7671 1000 7682 1034
rect 7626 966 7682 1000
rect 7626 932 7637 966
rect 7671 932 7682 966
rect 7626 898 7682 932
rect 7626 864 7637 898
rect 7671 864 7682 898
rect 7626 840 7682 864
rect 7712 1034 7768 1050
rect 7712 1000 7723 1034
rect 7757 1000 7768 1034
rect 7712 966 7768 1000
rect 7712 932 7723 966
rect 7757 932 7768 966
rect 7712 898 7768 932
rect 7712 864 7723 898
rect 7757 864 7768 898
rect 7712 840 7768 864
rect 7798 1034 7854 1050
rect 7798 1000 7809 1034
rect 7843 1000 7854 1034
rect 7798 966 7854 1000
rect 7798 932 7809 966
rect 7843 932 7854 966
rect 7798 898 7854 932
rect 7798 864 7809 898
rect 7843 864 7854 898
rect 7798 840 7854 864
rect 7884 1034 7940 1050
rect 7884 1000 7895 1034
rect 7929 1000 7940 1034
rect 7884 966 7940 1000
rect 7884 932 7895 966
rect 7929 932 7940 966
rect 7884 898 7940 932
rect 7884 864 7895 898
rect 7929 864 7940 898
rect 7884 840 7940 864
rect 7970 1034 8026 1050
rect 7970 1000 7981 1034
rect 8015 1000 8026 1034
rect 7970 966 8026 1000
rect 7970 932 7981 966
rect 8015 932 8026 966
rect 7970 898 8026 932
rect 7970 864 7981 898
rect 8015 864 8026 898
rect 7970 840 8026 864
rect 8056 1034 8112 1050
rect 8056 1000 8067 1034
rect 8101 1000 8112 1034
rect 8056 966 8112 1000
rect 8056 932 8067 966
rect 8101 932 8112 966
rect 8056 898 8112 932
rect 8056 864 8067 898
rect 8101 864 8112 898
rect 8056 840 8112 864
rect 8142 1034 8198 1050
rect 8142 1000 8153 1034
rect 8187 1000 8198 1034
rect 8142 966 8198 1000
rect 8142 932 8153 966
rect 8187 932 8198 966
rect 8142 898 8198 932
rect 8142 864 8153 898
rect 8187 864 8198 898
rect 8142 840 8198 864
rect 8228 1034 8284 1050
rect 8228 1000 8239 1034
rect 8273 1000 8284 1034
rect 8228 966 8284 1000
rect 8228 932 8239 966
rect 8273 932 8284 966
rect 8228 898 8284 932
rect 8228 864 8239 898
rect 8273 864 8284 898
rect 8228 840 8284 864
rect 8314 1034 8370 1050
rect 8314 1000 8325 1034
rect 8359 1000 8370 1034
rect 8314 966 8370 1000
rect 8314 932 8325 966
rect 8359 932 8370 966
rect 8314 898 8370 932
rect 8314 864 8325 898
rect 8359 864 8370 898
rect 8314 840 8370 864
rect 8400 1034 8456 1050
rect 8400 1000 8411 1034
rect 8445 1000 8456 1034
rect 8400 966 8456 1000
rect 8400 932 8411 966
rect 8445 932 8456 966
rect 8400 898 8456 932
rect 8400 864 8411 898
rect 8445 864 8456 898
rect 8400 840 8456 864
rect 8486 1034 8542 1050
rect 8486 1000 8497 1034
rect 8531 1000 8542 1034
rect 8486 966 8542 1000
rect 8486 932 8497 966
rect 8531 932 8542 966
rect 8486 898 8542 932
rect 8486 864 8497 898
rect 8531 864 8542 898
rect 8486 840 8542 864
rect 8572 1034 8628 1050
rect 8572 1000 8583 1034
rect 8617 1000 8628 1034
rect 8572 966 8628 1000
rect 8572 932 8583 966
rect 8617 932 8628 966
rect 8572 898 8628 932
rect 8572 864 8583 898
rect 8617 864 8628 898
rect 8572 840 8628 864
rect 8658 1034 8714 1050
rect 8658 1000 8669 1034
rect 8703 1000 8714 1034
rect 8658 966 8714 1000
rect 8658 932 8669 966
rect 8703 932 8714 966
rect 8658 898 8714 932
rect 8658 864 8669 898
rect 8703 864 8714 898
rect 8658 840 8714 864
rect 8744 1034 8800 1050
rect 8744 1000 8755 1034
rect 8789 1000 8800 1034
rect 8744 966 8800 1000
rect 8744 932 8755 966
rect 8789 932 8800 966
rect 8744 898 8800 932
rect 8744 864 8755 898
rect 8789 864 8800 898
rect 8744 840 8800 864
rect 8830 1034 8886 1050
rect 8830 1000 8841 1034
rect 8875 1000 8886 1034
rect 8830 966 8886 1000
rect 8830 932 8841 966
rect 8875 932 8886 966
rect 8830 898 8886 932
rect 8830 864 8841 898
rect 8875 864 8886 898
rect 8830 840 8886 864
rect 8916 1034 8972 1050
rect 8916 1000 8927 1034
rect 8961 1000 8972 1034
rect 8916 966 8972 1000
rect 8916 932 8927 966
rect 8961 932 8972 966
rect 8916 898 8972 932
rect 8916 864 8927 898
rect 8961 864 8972 898
rect 8916 840 8972 864
rect 9002 1034 9058 1050
rect 9002 1000 9013 1034
rect 9047 1000 9058 1034
rect 9002 966 9058 1000
rect 9002 932 9013 966
rect 9047 932 9058 966
rect 9002 898 9058 932
rect 9002 864 9013 898
rect 9047 864 9058 898
rect 9002 840 9058 864
rect 9088 1034 9144 1050
rect 9088 1000 9099 1034
rect 9133 1000 9144 1034
rect 9088 966 9144 1000
rect 9088 932 9099 966
rect 9133 932 9144 966
rect 9088 898 9144 932
rect 9088 864 9099 898
rect 9133 864 9144 898
rect 9088 840 9144 864
rect 9174 1034 9230 1050
rect 9174 1000 9185 1034
rect 9219 1000 9230 1034
rect 9174 966 9230 1000
rect 9174 932 9185 966
rect 9219 932 9230 966
rect 9174 898 9230 932
rect 9174 864 9185 898
rect 9219 864 9230 898
rect 9174 840 9230 864
rect 9260 1034 9316 1050
rect 9260 1000 9271 1034
rect 9305 1000 9316 1034
rect 9260 966 9316 1000
rect 9260 932 9271 966
rect 9305 932 9316 966
rect 9260 898 9316 932
rect 9260 864 9271 898
rect 9305 864 9316 898
rect 9260 840 9316 864
rect 9346 1034 9402 1050
rect 9346 1000 9357 1034
rect 9391 1000 9402 1034
rect 9346 966 9402 1000
rect 9346 932 9357 966
rect 9391 932 9402 966
rect 9346 898 9402 932
rect 9346 864 9357 898
rect 9391 864 9402 898
rect 9346 840 9402 864
rect 9432 1034 9488 1050
rect 9432 1000 9443 1034
rect 9477 1000 9488 1034
rect 9432 966 9488 1000
rect 9432 932 9443 966
rect 9477 932 9488 966
rect 9432 898 9488 932
rect 9432 864 9443 898
rect 9477 864 9488 898
rect 9432 840 9488 864
rect 9518 1034 9574 1050
rect 9518 1000 9529 1034
rect 9563 1000 9574 1034
rect 9518 966 9574 1000
rect 9518 932 9529 966
rect 9563 932 9574 966
rect 9518 898 9574 932
rect 9518 864 9529 898
rect 9563 864 9574 898
rect 9518 840 9574 864
rect 9604 1034 9660 1050
rect 9604 1000 9615 1034
rect 9649 1000 9660 1034
rect 9604 966 9660 1000
rect 9604 932 9615 966
rect 9649 932 9660 966
rect 9604 898 9660 932
rect 9604 864 9615 898
rect 9649 864 9660 898
rect 9604 840 9660 864
rect 9690 1034 9746 1050
rect 9690 1000 9701 1034
rect 9735 1000 9746 1034
rect 9690 966 9746 1000
rect 9690 932 9701 966
rect 9735 932 9746 966
rect 9690 898 9746 932
rect 9690 864 9701 898
rect 9735 864 9746 898
rect 9690 840 9746 864
rect 9776 1034 9832 1050
rect 9776 1000 9787 1034
rect 9821 1000 9832 1034
rect 9776 966 9832 1000
rect 9776 932 9787 966
rect 9821 932 9832 966
rect 9776 898 9832 932
rect 9776 864 9787 898
rect 9821 864 9832 898
rect 9776 840 9832 864
rect 9862 1034 9918 1050
rect 9862 1000 9873 1034
rect 9907 1000 9918 1034
rect 9862 966 9918 1000
rect 9862 932 9873 966
rect 9907 932 9918 966
rect 9862 898 9918 932
rect 9862 864 9873 898
rect 9907 864 9918 898
rect 9862 840 9918 864
rect 9948 1034 10004 1050
rect 9948 1000 9959 1034
rect 9993 1000 10004 1034
rect 9948 966 10004 1000
rect 9948 932 9959 966
rect 9993 932 10004 966
rect 9948 898 10004 932
rect 9948 864 9959 898
rect 9993 864 10004 898
rect 9948 840 10004 864
rect 10034 1034 10090 1050
rect 10034 1000 10045 1034
rect 10079 1000 10090 1034
rect 10034 966 10090 1000
rect 10034 932 10045 966
rect 10079 932 10090 966
rect 10034 898 10090 932
rect 10034 864 10045 898
rect 10079 864 10090 898
rect 10034 840 10090 864
rect 10120 1034 10176 1050
rect 10120 1000 10131 1034
rect 10165 1000 10176 1034
rect 10120 966 10176 1000
rect 10120 932 10131 966
rect 10165 932 10176 966
rect 10120 898 10176 932
rect 10120 864 10131 898
rect 10165 864 10176 898
rect 10120 840 10176 864
rect 10206 1034 10262 1050
rect 10206 1000 10217 1034
rect 10251 1000 10262 1034
rect 10206 966 10262 1000
rect 10206 932 10217 966
rect 10251 932 10262 966
rect 10206 898 10262 932
rect 10206 864 10217 898
rect 10251 864 10262 898
rect 10206 840 10262 864
rect 10292 1034 10348 1050
rect 10292 1000 10303 1034
rect 10337 1000 10348 1034
rect 10292 966 10348 1000
rect 10292 932 10303 966
rect 10337 932 10348 966
rect 10292 898 10348 932
rect 10292 864 10303 898
rect 10337 864 10348 898
rect 10292 840 10348 864
rect 10378 1034 10434 1050
rect 10378 1000 10389 1034
rect 10423 1000 10434 1034
rect 10378 966 10434 1000
rect 10378 932 10389 966
rect 10423 932 10434 966
rect 10378 898 10434 932
rect 10378 864 10389 898
rect 10423 864 10434 898
rect 10378 840 10434 864
rect 10464 1034 10520 1050
rect 10464 1000 10475 1034
rect 10509 1000 10520 1034
rect 10464 966 10520 1000
rect 10464 932 10475 966
rect 10509 932 10520 966
rect 10464 898 10520 932
rect 10464 864 10475 898
rect 10509 864 10520 898
rect 10464 840 10520 864
rect 10550 1034 10606 1050
rect 10550 1000 10561 1034
rect 10595 1000 10606 1034
rect 10550 966 10606 1000
rect 10550 932 10561 966
rect 10595 932 10606 966
rect 10550 898 10606 932
rect 10550 864 10561 898
rect 10595 864 10606 898
rect 10550 840 10606 864
rect 10636 1034 10692 1050
rect 10636 1000 10647 1034
rect 10681 1000 10692 1034
rect 10636 966 10692 1000
rect 10636 932 10647 966
rect 10681 932 10692 966
rect 10636 898 10692 932
rect 10636 864 10647 898
rect 10681 864 10692 898
rect 10636 840 10692 864
rect 10722 1034 10778 1050
rect 10722 1000 10733 1034
rect 10767 1000 10778 1034
rect 10722 966 10778 1000
rect 10722 932 10733 966
rect 10767 932 10778 966
rect 10722 898 10778 932
rect 10722 864 10733 898
rect 10767 864 10778 898
rect 10722 840 10778 864
rect 10808 1034 10864 1050
rect 10808 1000 10819 1034
rect 10853 1000 10864 1034
rect 10808 966 10864 1000
rect 10808 932 10819 966
rect 10853 932 10864 966
rect 10808 898 10864 932
rect 10808 864 10819 898
rect 10853 864 10864 898
rect 10808 840 10864 864
rect 10894 1034 10950 1050
rect 10894 1000 10905 1034
rect 10939 1000 10950 1034
rect 10894 966 10950 1000
rect 10894 932 10905 966
rect 10939 932 10950 966
rect 10894 898 10950 932
rect 10894 864 10905 898
rect 10939 864 10950 898
rect 10894 840 10950 864
rect 10980 1034 11036 1050
rect 10980 1000 10991 1034
rect 11025 1000 11036 1034
rect 10980 966 11036 1000
rect 10980 932 10991 966
rect 11025 932 11036 966
rect 10980 898 11036 932
rect 10980 864 10991 898
rect 11025 864 11036 898
rect 10980 840 11036 864
rect 11066 1034 11122 1050
rect 11066 1000 11077 1034
rect 11111 1000 11122 1034
rect 11066 966 11122 1000
rect 11066 932 11077 966
rect 11111 932 11122 966
rect 11066 898 11122 932
rect 11066 864 11077 898
rect 11111 864 11122 898
rect 11066 840 11122 864
rect 11152 1034 11208 1050
rect 11152 1000 11163 1034
rect 11197 1000 11208 1034
rect 11152 966 11208 1000
rect 11152 932 11163 966
rect 11197 932 11208 966
rect 11152 898 11208 932
rect 11152 864 11163 898
rect 11197 864 11208 898
rect 11152 840 11208 864
rect 11238 1034 11294 1050
rect 11238 1000 11249 1034
rect 11283 1000 11294 1034
rect 11238 966 11294 1000
rect 11238 932 11249 966
rect 11283 932 11294 966
rect 11238 898 11294 932
rect 11238 864 11249 898
rect 11283 864 11294 898
rect 11238 840 11294 864
rect 11324 1034 11377 1050
rect 11324 1000 11335 1034
rect 11369 1000 11377 1034
rect 11324 966 11377 1000
rect 11324 932 11335 966
rect 11369 932 11377 966
rect 11324 898 11377 932
rect 11324 864 11335 898
rect 11369 864 11377 898
rect 11324 840 11377 864
<< ndiffc >>
rect 1101 3302 1135 3336
rect 1101 3234 1135 3268
rect 1101 3166 1135 3200
rect 1187 3302 1221 3336
rect 1187 3234 1221 3268
rect 1187 3166 1221 3200
rect 1273 3302 1307 3336
rect 1273 3234 1307 3268
rect 1273 3166 1307 3200
rect 2993 3302 3027 3336
rect 2993 3234 3027 3268
rect 2993 3166 3027 3200
rect 3079 3302 3113 3336
rect 3079 3234 3113 3268
rect 3079 3166 3113 3200
rect 3165 3302 3199 3336
rect 3165 3234 3199 3268
rect 3165 3166 3199 3200
rect 6691 3302 6725 3336
rect 6691 3234 6725 3268
rect 6691 3166 6725 3200
rect 6777 3302 6811 3336
rect 6777 3234 6811 3268
rect 6777 3166 6811 3200
rect 6863 3302 6897 3336
rect 6863 3234 6897 3268
rect 6863 3166 6897 3200
rect 9185 3302 9219 3336
rect 9185 3234 9219 3268
rect 9185 3166 9219 3200
rect 9271 3302 9305 3336
rect 9271 3234 9305 3268
rect 9271 3166 9305 3200
rect 9357 3302 9391 3336
rect 9357 3234 9391 3268
rect 9357 3166 9391 3200
rect 6175 2966 6209 3000
rect 6175 2898 6209 2932
rect 6175 2830 6209 2864
rect 6261 2966 6295 3000
rect 6261 2898 6295 2932
rect 6261 2830 6295 2864
rect 6347 2966 6381 3000
rect 6347 2898 6381 2932
rect 6347 2830 6381 2864
rect 4369 2546 4403 2580
rect 4369 2478 4403 2512
rect 4369 2410 4403 2444
rect 4455 2546 4489 2580
rect 4455 2478 4489 2512
rect 4455 2410 4489 2444
rect 4541 2546 4575 2580
rect 4541 2478 4575 2512
rect 4541 2410 4575 2444
rect 5487 2546 5521 2580
rect 5487 2478 5521 2512
rect 5487 2410 5521 2444
rect 5573 2546 5607 2580
rect 5573 2478 5607 2512
rect 5573 2410 5607 2444
rect 5659 2546 5693 2580
rect 5659 2478 5693 2512
rect 5659 2410 5693 2444
rect 6175 1454 6209 1488
rect 6175 1386 6209 1420
rect 6175 1318 6209 1352
rect 6261 1454 6295 1488
rect 6261 1386 6295 1420
rect 6261 1318 6295 1352
rect 6347 1454 6381 1488
rect 6347 1386 6381 1420
rect 6347 1318 6381 1352
<< pdiffc >>
rect 155 2176 189 2210
rect 155 2108 189 2142
rect 155 2040 189 2074
rect 241 2176 275 2210
rect 241 2108 275 2142
rect 241 2040 275 2074
rect 327 2176 361 2210
rect 327 2108 361 2142
rect 327 2040 361 2074
rect 413 2176 447 2210
rect 413 2108 447 2142
rect 413 2040 447 2074
rect 499 2176 533 2210
rect 499 2108 533 2142
rect 499 2040 533 2074
rect 585 2176 619 2210
rect 585 2108 619 2142
rect 585 2040 619 2074
rect 671 2176 705 2210
rect 671 2108 705 2142
rect 671 2040 705 2074
rect 757 2176 791 2210
rect 757 2108 791 2142
rect 757 2040 791 2074
rect 843 2176 877 2210
rect 843 2108 877 2142
rect 843 2040 877 2074
rect 929 2176 963 2210
rect 929 2108 963 2142
rect 929 2040 963 2074
rect 1015 2176 1049 2210
rect 1015 2108 1049 2142
rect 1015 2040 1049 2074
rect 1101 2176 1135 2210
rect 1101 2108 1135 2142
rect 1101 2040 1135 2074
rect 1187 2176 1221 2210
rect 1187 2108 1221 2142
rect 1187 2040 1221 2074
rect 1273 2176 1307 2210
rect 1273 2108 1307 2142
rect 1273 2040 1307 2074
rect 1359 2176 1393 2210
rect 1359 2108 1393 2142
rect 1359 2040 1393 2074
rect 1445 2176 1479 2210
rect 1445 2108 1479 2142
rect 1445 2040 1479 2074
rect 1531 2176 1565 2210
rect 1531 2108 1565 2142
rect 1531 2040 1565 2074
rect 1617 2176 1651 2210
rect 1617 2108 1651 2142
rect 1617 2040 1651 2074
rect 1703 2176 1737 2210
rect 1703 2108 1737 2142
rect 1703 2040 1737 2074
rect 1789 2176 1823 2210
rect 1789 2108 1823 2142
rect 1789 2040 1823 2074
rect 1875 2176 1909 2210
rect 1875 2108 1909 2142
rect 1875 2040 1909 2074
rect 1961 2176 1995 2210
rect 1961 2108 1995 2142
rect 1961 2040 1995 2074
rect 2047 2176 2081 2210
rect 2047 2108 2081 2142
rect 2047 2040 2081 2074
rect 2133 2176 2167 2210
rect 2133 2108 2167 2142
rect 2133 2040 2167 2074
rect 2219 2176 2253 2210
rect 2219 2108 2253 2142
rect 2219 2040 2253 2074
rect 2563 2176 2597 2210
rect 2563 2108 2597 2142
rect 2563 2040 2597 2074
rect 2649 2176 2683 2210
rect 2649 2108 2683 2142
rect 2649 2040 2683 2074
rect 2735 2176 2769 2210
rect 2735 2108 2769 2142
rect 2735 2040 2769 2074
rect 2821 2176 2855 2210
rect 2821 2108 2855 2142
rect 2821 2040 2855 2074
rect 2907 2176 2941 2210
rect 2907 2108 2941 2142
rect 2907 2040 2941 2074
rect 2993 2176 3027 2210
rect 2993 2108 3027 2142
rect 2993 2040 3027 2074
rect 3079 2176 3113 2210
rect 3079 2108 3113 2142
rect 3079 2040 3113 2074
rect 3165 2176 3199 2210
rect 3165 2108 3199 2142
rect 3165 2040 3199 2074
rect 3251 2176 3285 2210
rect 3251 2108 3285 2142
rect 3251 2040 3285 2074
rect 3337 2176 3371 2210
rect 3337 2108 3371 2142
rect 3337 2040 3371 2074
rect 3423 2176 3457 2210
rect 3423 2108 3457 2142
rect 3423 2040 3457 2074
rect 3509 2176 3543 2210
rect 3509 2108 3543 2142
rect 3509 2040 3543 2074
rect 3595 2176 3629 2210
rect 3595 2108 3629 2142
rect 3595 2040 3629 2074
rect 6691 2176 6725 2210
rect 6691 2108 6725 2142
rect 6691 2040 6725 2074
rect 6777 2176 6811 2210
rect 6777 2108 6811 2142
rect 6777 2040 6811 2074
rect 6863 2176 6897 2210
rect 6863 2108 6897 2142
rect 6863 2040 6897 2074
rect 7207 2176 7241 2210
rect 7207 2108 7241 2142
rect 7207 2040 7241 2074
rect 7293 2176 7327 2210
rect 7293 2108 7327 2142
rect 7293 2040 7327 2074
rect 7379 2176 7413 2210
rect 7379 2108 7413 2142
rect 7379 2040 7413 2074
rect 7465 2176 7499 2210
rect 7465 2108 7499 2142
rect 7465 2040 7499 2074
rect 7551 2176 7585 2210
rect 7551 2108 7585 2142
rect 7551 2040 7585 2074
rect 7637 2176 7671 2210
rect 7637 2108 7671 2142
rect 7637 2040 7671 2074
rect 7723 2176 7757 2210
rect 7723 2108 7757 2142
rect 7723 2040 7757 2074
rect 7809 2176 7843 2210
rect 7809 2108 7843 2142
rect 7809 2040 7843 2074
rect 7895 2176 7929 2210
rect 7895 2108 7929 2142
rect 7895 2040 7929 2074
rect 7981 2176 8015 2210
rect 7981 2108 8015 2142
rect 7981 2040 8015 2074
rect 8067 2176 8101 2210
rect 8067 2108 8101 2142
rect 8067 2040 8101 2074
rect 8153 2176 8187 2210
rect 8153 2108 8187 2142
rect 8153 2040 8187 2074
rect 8239 2176 8273 2210
rect 8239 2108 8273 2142
rect 8239 2040 8273 2074
rect 8325 2176 8359 2210
rect 8325 2108 8359 2142
rect 8325 2040 8359 2074
rect 8411 2176 8445 2210
rect 8411 2108 8445 2142
rect 8411 2040 8445 2074
rect 8497 2176 8531 2210
rect 8497 2108 8531 2142
rect 8497 2040 8531 2074
rect 8583 2176 8617 2210
rect 8583 2108 8617 2142
rect 8583 2040 8617 2074
rect 8669 2176 8703 2210
rect 8669 2108 8703 2142
rect 8669 2040 8703 2074
rect 8755 2176 8789 2210
rect 8755 2108 8789 2142
rect 8755 2040 8789 2074
rect 8841 2176 8875 2210
rect 8841 2108 8875 2142
rect 8841 2040 8875 2074
rect 8927 2176 8961 2210
rect 8927 2108 8961 2142
rect 8927 2040 8961 2074
rect 9013 2176 9047 2210
rect 9013 2108 9047 2142
rect 9013 2040 9047 2074
rect 9099 2176 9133 2210
rect 9099 2108 9133 2142
rect 9099 2040 9133 2074
rect 9185 2176 9219 2210
rect 9185 2108 9219 2142
rect 9185 2040 9219 2074
rect 9271 2176 9305 2210
rect 9271 2108 9305 2142
rect 9271 2040 9305 2074
rect 9357 2176 9391 2210
rect 9357 2108 9391 2142
rect 9357 2040 9391 2074
rect 9443 2176 9477 2210
rect 9443 2108 9477 2142
rect 9443 2040 9477 2074
rect 9529 2176 9563 2210
rect 9529 2108 9563 2142
rect 9529 2040 9563 2074
rect 9615 2176 9649 2210
rect 9615 2108 9649 2142
rect 9615 2040 9649 2074
rect 9701 2176 9735 2210
rect 9701 2108 9735 2142
rect 9701 2040 9735 2074
rect 9787 2176 9821 2210
rect 9787 2108 9821 2142
rect 9787 2040 9821 2074
rect 9873 2176 9907 2210
rect 9873 2108 9907 2142
rect 9873 2040 9907 2074
rect 9959 2176 9993 2210
rect 9959 2108 9993 2142
rect 9959 2040 9993 2074
rect 10045 2176 10079 2210
rect 10045 2108 10079 2142
rect 10045 2040 10079 2074
rect 10131 2176 10165 2210
rect 10131 2108 10165 2142
rect 10131 2040 10165 2074
rect 10217 2176 10251 2210
rect 10217 2108 10251 2142
rect 10217 2040 10251 2074
rect 10303 2176 10337 2210
rect 10303 2108 10337 2142
rect 10303 2040 10337 2074
rect 10389 2176 10423 2210
rect 10389 2108 10423 2142
rect 10389 2040 10423 2074
rect 10475 2176 10509 2210
rect 10475 2108 10509 2142
rect 10475 2040 10509 2074
rect 10561 2176 10595 2210
rect 10561 2108 10595 2142
rect 10561 2040 10595 2074
rect 10647 2176 10681 2210
rect 10647 2108 10681 2142
rect 10647 2040 10681 2074
rect 10733 2176 10767 2210
rect 10733 2108 10767 2142
rect 10733 2040 10767 2074
rect 10819 2176 10853 2210
rect 10819 2108 10853 2142
rect 10819 2040 10853 2074
rect 10905 2176 10939 2210
rect 10905 2108 10939 2142
rect 10905 2040 10939 2074
rect 10991 2176 11025 2210
rect 10991 2108 11025 2142
rect 10991 2040 11025 2074
rect 11077 2176 11111 2210
rect 11077 2108 11111 2142
rect 11077 2040 11111 2074
rect 11163 2176 11197 2210
rect 11163 2108 11197 2142
rect 11163 2040 11197 2074
rect 11249 2176 11283 2210
rect 11249 2108 11283 2142
rect 11249 2040 11283 2074
rect 11335 2176 11369 2210
rect 11335 2108 11369 2142
rect 11335 2040 11369 2074
rect 3939 1420 3973 1454
rect 3939 1352 3973 1386
rect 3939 1284 3973 1318
rect 4025 1420 4059 1454
rect 4025 1352 4059 1386
rect 4025 1284 4059 1318
rect 4111 1420 4145 1454
rect 4111 1352 4145 1386
rect 4111 1284 4145 1318
rect 4197 1420 4231 1454
rect 4197 1352 4231 1386
rect 4197 1284 4231 1318
rect 4283 1420 4317 1454
rect 4283 1352 4317 1386
rect 4283 1284 4317 1318
rect 4369 1420 4403 1454
rect 4369 1352 4403 1386
rect 4369 1284 4403 1318
rect 4455 1420 4489 1454
rect 4455 1352 4489 1386
rect 4455 1284 4489 1318
rect 4541 1420 4575 1454
rect 4541 1352 4575 1386
rect 4541 1284 4575 1318
rect 4627 1420 4661 1454
rect 4627 1352 4661 1386
rect 4627 1284 4661 1318
rect 4713 1420 4747 1454
rect 4713 1352 4747 1386
rect 4713 1284 4747 1318
rect 4799 1420 4833 1454
rect 4799 1352 4833 1386
rect 4799 1284 4833 1318
rect 4885 1420 4919 1454
rect 4885 1352 4919 1386
rect 4885 1284 4919 1318
rect 4971 1420 5005 1454
rect 4971 1352 5005 1386
rect 4971 1284 5005 1318
rect 5315 1420 5349 1454
rect 5315 1352 5349 1386
rect 5315 1284 5349 1318
rect 5401 1420 5435 1454
rect 5401 1352 5435 1386
rect 5401 1284 5435 1318
rect 5487 1420 5521 1454
rect 5487 1352 5521 1386
rect 5487 1284 5521 1318
rect 5573 1420 5607 1454
rect 5573 1352 5607 1386
rect 5573 1284 5607 1318
rect 5659 1420 5693 1454
rect 5659 1352 5693 1386
rect 5659 1284 5693 1318
rect 5745 1420 5779 1454
rect 5745 1352 5779 1386
rect 5745 1284 5779 1318
rect 5831 1420 5865 1454
rect 5831 1352 5865 1386
rect 5831 1284 5865 1318
rect 155 1000 189 1034
rect 155 932 189 966
rect 155 864 189 898
rect 241 1000 275 1034
rect 241 932 275 966
rect 241 864 275 898
rect 327 1000 361 1034
rect 327 932 361 966
rect 327 864 361 898
rect 413 1000 447 1034
rect 413 932 447 966
rect 413 864 447 898
rect 499 1000 533 1034
rect 499 932 533 966
rect 499 864 533 898
rect 585 1000 619 1034
rect 585 932 619 966
rect 585 864 619 898
rect 671 1000 705 1034
rect 671 932 705 966
rect 671 864 705 898
rect 757 1000 791 1034
rect 757 932 791 966
rect 757 864 791 898
rect 843 1000 877 1034
rect 843 932 877 966
rect 843 864 877 898
rect 929 1000 963 1034
rect 929 932 963 966
rect 929 864 963 898
rect 1015 1000 1049 1034
rect 1015 932 1049 966
rect 1015 864 1049 898
rect 1101 1000 1135 1034
rect 1101 932 1135 966
rect 1101 864 1135 898
rect 1187 1000 1221 1034
rect 1187 932 1221 966
rect 1187 864 1221 898
rect 1273 1000 1307 1034
rect 1273 932 1307 966
rect 1273 864 1307 898
rect 1359 1000 1393 1034
rect 1359 932 1393 966
rect 1359 864 1393 898
rect 1445 1000 1479 1034
rect 1445 932 1479 966
rect 1445 864 1479 898
rect 1531 1000 1565 1034
rect 1531 932 1565 966
rect 1531 864 1565 898
rect 1617 1000 1651 1034
rect 1617 932 1651 966
rect 1617 864 1651 898
rect 1703 1000 1737 1034
rect 1703 932 1737 966
rect 1703 864 1737 898
rect 1789 1000 1823 1034
rect 1789 932 1823 966
rect 1789 864 1823 898
rect 1875 1000 1909 1034
rect 1875 932 1909 966
rect 1875 864 1909 898
rect 1961 1000 1995 1034
rect 1961 932 1995 966
rect 1961 864 1995 898
rect 2047 1000 2081 1034
rect 2047 932 2081 966
rect 2047 864 2081 898
rect 2133 1000 2167 1034
rect 2133 932 2167 966
rect 2133 864 2167 898
rect 2219 1000 2253 1034
rect 2219 932 2253 966
rect 2219 864 2253 898
rect 2563 1000 2597 1034
rect 2563 932 2597 966
rect 2563 864 2597 898
rect 2649 1000 2683 1034
rect 2649 932 2683 966
rect 2649 864 2683 898
rect 2735 1000 2769 1034
rect 2735 932 2769 966
rect 2735 864 2769 898
rect 2821 1000 2855 1034
rect 2821 932 2855 966
rect 2821 864 2855 898
rect 2907 1000 2941 1034
rect 2907 932 2941 966
rect 2907 864 2941 898
rect 2993 1000 3027 1034
rect 2993 932 3027 966
rect 2993 864 3027 898
rect 3079 1000 3113 1034
rect 3079 932 3113 966
rect 3079 864 3113 898
rect 3165 1000 3199 1034
rect 3165 932 3199 966
rect 3165 864 3199 898
rect 3251 1000 3285 1034
rect 3251 932 3285 966
rect 3251 864 3285 898
rect 3337 1000 3371 1034
rect 3337 932 3371 966
rect 3337 864 3371 898
rect 3423 1000 3457 1034
rect 3423 932 3457 966
rect 3423 864 3457 898
rect 3509 1000 3543 1034
rect 3509 932 3543 966
rect 3509 864 3543 898
rect 3595 1000 3629 1034
rect 7207 1000 7241 1034
rect 3595 932 3629 966
rect 3595 864 3629 898
rect 7207 932 7241 966
rect 7207 864 7241 898
rect 7293 1000 7327 1034
rect 7293 932 7327 966
rect 7293 864 7327 898
rect 7379 1000 7413 1034
rect 7379 932 7413 966
rect 7379 864 7413 898
rect 7465 1000 7499 1034
rect 7465 932 7499 966
rect 7465 864 7499 898
rect 7551 1000 7585 1034
rect 7551 932 7585 966
rect 7551 864 7585 898
rect 7637 1000 7671 1034
rect 7637 932 7671 966
rect 7637 864 7671 898
rect 7723 1000 7757 1034
rect 7723 932 7757 966
rect 7723 864 7757 898
rect 7809 1000 7843 1034
rect 7809 932 7843 966
rect 7809 864 7843 898
rect 7895 1000 7929 1034
rect 7895 932 7929 966
rect 7895 864 7929 898
rect 7981 1000 8015 1034
rect 7981 932 8015 966
rect 7981 864 8015 898
rect 8067 1000 8101 1034
rect 8067 932 8101 966
rect 8067 864 8101 898
rect 8153 1000 8187 1034
rect 8153 932 8187 966
rect 8153 864 8187 898
rect 8239 1000 8273 1034
rect 8239 932 8273 966
rect 8239 864 8273 898
rect 8325 1000 8359 1034
rect 8325 932 8359 966
rect 8325 864 8359 898
rect 8411 1000 8445 1034
rect 8411 932 8445 966
rect 8411 864 8445 898
rect 8497 1000 8531 1034
rect 8497 932 8531 966
rect 8497 864 8531 898
rect 8583 1000 8617 1034
rect 8583 932 8617 966
rect 8583 864 8617 898
rect 8669 1000 8703 1034
rect 8669 932 8703 966
rect 8669 864 8703 898
rect 8755 1000 8789 1034
rect 8755 932 8789 966
rect 8755 864 8789 898
rect 8841 1000 8875 1034
rect 8841 932 8875 966
rect 8841 864 8875 898
rect 8927 1000 8961 1034
rect 8927 932 8961 966
rect 8927 864 8961 898
rect 9013 1000 9047 1034
rect 9013 932 9047 966
rect 9013 864 9047 898
rect 9099 1000 9133 1034
rect 9099 932 9133 966
rect 9099 864 9133 898
rect 9185 1000 9219 1034
rect 9185 932 9219 966
rect 9185 864 9219 898
rect 9271 1000 9305 1034
rect 9271 932 9305 966
rect 9271 864 9305 898
rect 9357 1000 9391 1034
rect 9357 932 9391 966
rect 9357 864 9391 898
rect 9443 1000 9477 1034
rect 9443 932 9477 966
rect 9443 864 9477 898
rect 9529 1000 9563 1034
rect 9529 932 9563 966
rect 9529 864 9563 898
rect 9615 1000 9649 1034
rect 9615 932 9649 966
rect 9615 864 9649 898
rect 9701 1000 9735 1034
rect 9701 932 9735 966
rect 9701 864 9735 898
rect 9787 1000 9821 1034
rect 9787 932 9821 966
rect 9787 864 9821 898
rect 9873 1000 9907 1034
rect 9873 932 9907 966
rect 9873 864 9907 898
rect 9959 1000 9993 1034
rect 9959 932 9993 966
rect 9959 864 9993 898
rect 10045 1000 10079 1034
rect 10045 932 10079 966
rect 10045 864 10079 898
rect 10131 1000 10165 1034
rect 10131 932 10165 966
rect 10131 864 10165 898
rect 10217 1000 10251 1034
rect 10217 932 10251 966
rect 10217 864 10251 898
rect 10303 1000 10337 1034
rect 10303 932 10337 966
rect 10303 864 10337 898
rect 10389 1000 10423 1034
rect 10389 932 10423 966
rect 10389 864 10423 898
rect 10475 1000 10509 1034
rect 10475 932 10509 966
rect 10475 864 10509 898
rect 10561 1000 10595 1034
rect 10561 932 10595 966
rect 10561 864 10595 898
rect 10647 1000 10681 1034
rect 10647 932 10681 966
rect 10647 864 10681 898
rect 10733 1000 10767 1034
rect 10733 932 10767 966
rect 10733 864 10767 898
rect 10819 1000 10853 1034
rect 10819 932 10853 966
rect 10819 864 10853 898
rect 10905 1000 10939 1034
rect 10905 932 10939 966
rect 10905 864 10939 898
rect 10991 1000 11025 1034
rect 10991 932 11025 966
rect 10991 864 11025 898
rect 11077 1000 11111 1034
rect 11077 932 11111 966
rect 11077 864 11111 898
rect 11163 1000 11197 1034
rect 11163 932 11197 966
rect 11163 864 11197 898
rect 11249 1000 11283 1034
rect 11249 932 11283 966
rect 11249 864 11283 898
rect 11335 1000 11369 1034
rect 11335 932 11369 966
rect 11335 864 11369 898
<< psubdiff >>
rect 1187 4049 1221 4144
rect 1187 3920 1221 4015
rect 3079 4049 3113 4144
rect 3079 3920 3113 4015
rect 6777 4049 6811 4144
rect 6777 3920 6811 4015
rect 9271 4049 9305 4144
rect 9271 3920 9305 4015
rect 6261 3713 6295 3808
rect 6261 3584 6295 3679
rect 4455 3293 4489 3388
rect 4455 3164 4489 3259
rect 5573 3293 5607 3388
rect 5573 3164 5607 3259
rect 6261 2201 6295 2296
rect 6261 2072 6295 2167
<< nsubdiff >>
rect 6777 1361 6811 1456
rect 6777 1232 6811 1327
rect 4025 605 4059 700
rect 4025 476 4059 571
rect 4197 605 4231 700
rect 4197 476 4231 571
rect 4369 605 4403 700
rect 4369 476 4403 571
rect 4541 605 4575 700
rect 4541 476 4575 571
rect 4713 605 4747 700
rect 4713 476 4747 571
rect 4885 605 4919 700
rect 4885 476 4919 571
rect 5401 605 5435 700
rect 5401 476 5435 571
rect 5573 605 5607 700
rect 5573 476 5607 571
rect 5745 605 5779 700
rect 5745 476 5779 571
rect 241 185 275 280
rect 241 56 275 151
rect 413 185 447 280
rect 413 56 447 151
rect 585 185 619 280
rect 585 56 619 151
rect 757 185 791 280
rect 757 56 791 151
rect 929 185 963 280
rect 929 56 963 151
rect 1101 185 1135 280
rect 1101 56 1135 151
rect 1273 185 1307 280
rect 1273 56 1307 151
rect 1445 185 1479 280
rect 1445 56 1479 151
rect 1617 185 1651 280
rect 1617 56 1651 151
rect 1789 185 1823 280
rect 1789 56 1823 151
rect 1961 185 1995 280
rect 1961 56 1995 151
rect 2133 185 2167 280
rect 2133 56 2167 151
rect 2649 185 2683 280
rect 2649 56 2683 151
rect 2821 185 2855 280
rect 2821 56 2855 151
rect 2993 185 3027 280
rect 2993 56 3027 151
rect 3165 185 3199 280
rect 3165 56 3199 151
rect 3337 185 3371 280
rect 3337 56 3371 151
rect 3509 185 3543 280
rect 3509 56 3543 151
rect 7293 185 7327 280
rect 7293 56 7327 151
rect 7465 185 7499 280
rect 7465 56 7499 151
rect 7637 185 7671 280
rect 7637 56 7671 151
rect 7809 185 7843 280
rect 7809 56 7843 151
rect 7981 185 8015 280
rect 7981 56 8015 151
rect 8153 185 8187 280
rect 8153 56 8187 151
rect 8325 185 8359 280
rect 8325 56 8359 151
rect 8497 185 8531 280
rect 8497 56 8531 151
rect 8669 185 8703 280
rect 8669 56 8703 151
rect 8841 185 8875 280
rect 8841 56 8875 151
rect 9013 185 9047 280
rect 9013 56 9047 151
rect 9185 185 9219 280
rect 9185 56 9219 151
rect 9357 185 9391 280
rect 9357 56 9391 151
rect 9529 185 9563 280
rect 9529 56 9563 151
rect 9701 185 9735 280
rect 9701 56 9735 151
rect 9873 185 9907 280
rect 9873 56 9907 151
rect 10045 185 10079 280
rect 10045 56 10079 151
rect 10217 185 10251 280
rect 10217 56 10251 151
rect 10389 185 10423 280
rect 10389 56 10423 151
rect 10561 185 10595 280
rect 10561 56 10595 151
rect 10733 185 10767 280
rect 10733 56 10767 151
rect 10905 185 10939 280
rect 10905 56 10939 151
rect 11077 185 11111 280
rect 11077 56 11111 151
rect 11249 185 11283 280
rect 11249 56 11283 151
<< psubdiffcont >>
rect 1187 4015 1221 4049
rect 3079 4015 3113 4049
rect 6777 4015 6811 4049
rect 9271 4015 9305 4049
rect 6261 3679 6295 3713
rect 4455 3259 4489 3293
rect 5573 3259 5607 3293
rect 6261 2167 6295 2201
<< nsubdiffcont >>
rect 6777 1327 6811 1361
rect 4025 571 4059 605
rect 4197 571 4231 605
rect 4369 571 4403 605
rect 4541 571 4575 605
rect 4713 571 4747 605
rect 4885 571 4919 605
rect 5401 571 5435 605
rect 5573 571 5607 605
rect 5745 571 5779 605
rect 241 151 275 185
rect 413 151 447 185
rect 585 151 619 185
rect 757 151 791 185
rect 929 151 963 185
rect 1101 151 1135 185
rect 1273 151 1307 185
rect 1445 151 1479 185
rect 1617 151 1651 185
rect 1789 151 1823 185
rect 1961 151 1995 185
rect 2133 151 2167 185
rect 2649 151 2683 185
rect 2821 151 2855 185
rect 2993 151 3027 185
rect 3165 151 3199 185
rect 3337 151 3371 185
rect 3509 151 3543 185
rect 7293 151 7327 185
rect 7465 151 7499 185
rect 7637 151 7671 185
rect 7809 151 7843 185
rect 7981 151 8015 185
rect 8153 151 8187 185
rect 8325 151 8359 185
rect 8497 151 8531 185
rect 8669 151 8703 185
rect 8841 151 8875 185
rect 9013 151 9047 185
rect 9185 151 9219 185
rect 9357 151 9391 185
rect 9529 151 9563 185
rect 9701 151 9735 185
rect 9873 151 9907 185
rect 10045 151 10079 185
rect 10217 151 10251 185
rect 10389 151 10423 185
rect 10561 151 10595 185
rect 10733 151 10767 185
rect 10905 151 10939 185
rect 11077 151 11111 185
rect 11249 151 11283 185
<< poly >>
rect 1146 3629 1262 3639
rect 1146 3595 1187 3629
rect 1221 3595 1262 3629
rect 1146 3585 1262 3595
rect 1146 3360 1176 3585
rect 1232 3360 1262 3585
rect 3038 3629 3154 3639
rect 3038 3595 3079 3629
rect 3113 3595 3154 3629
rect 3038 3585 3154 3595
rect 3038 3360 3068 3585
rect 3124 3360 3154 3585
rect 6736 3629 6852 3639
rect 6736 3595 6777 3629
rect 6811 3595 6852 3629
rect 6736 3585 6852 3595
rect 6736 3360 6766 3585
rect 6822 3360 6852 3585
rect 9230 3629 9346 3639
rect 9230 3595 9271 3629
rect 9305 3595 9346 3629
rect 9230 3585 9346 3595
rect 9230 3360 9260 3585
rect 9316 3360 9346 3585
rect 6220 3293 6336 3303
rect 6220 3259 6261 3293
rect 6295 3259 6336 3293
rect 6220 3249 6336 3259
rect 1146 2940 1176 3150
rect 1232 2940 1262 3150
rect 3038 2940 3068 3150
rect 3124 2940 3154 3150
rect 6220 3024 6250 3249
rect 6306 3024 6336 3249
rect 4414 2873 4530 2883
rect 4414 2839 4455 2873
rect 4489 2839 4530 2873
rect 4414 2829 4530 2839
rect 4414 2604 4444 2829
rect 4500 2604 4530 2829
rect 5532 2873 5648 2883
rect 5532 2839 5573 2873
rect 5607 2839 5648 2873
rect 5532 2829 5648 2839
rect 5532 2604 5562 2829
rect 5618 2604 5648 2829
rect 6736 2940 6766 3150
rect 6822 2940 6852 3150
rect 9230 2940 9260 3150
rect 9316 2940 9346 3150
rect 6220 2604 6250 2814
rect 6306 2604 6336 2814
rect 200 2226 230 2436
rect 286 2226 316 2436
rect 372 2226 402 2436
rect 458 2226 488 2436
rect 544 2226 574 2436
rect 630 2226 660 2436
rect 716 2226 746 2436
rect 802 2226 832 2436
rect 888 2226 918 2436
rect 974 2226 1004 2436
rect 1060 2226 1090 2436
rect 1146 2226 1176 2436
rect 1232 2226 1262 2436
rect 1318 2226 1348 2436
rect 1404 2226 1434 2436
rect 1490 2226 1520 2436
rect 1576 2226 1606 2436
rect 1662 2226 1692 2436
rect 1748 2226 1778 2436
rect 1834 2226 1864 2436
rect 1920 2226 1950 2436
rect 2006 2226 2036 2436
rect 2092 2226 2122 2436
rect 2178 2226 2208 2436
rect 2608 2226 2638 2436
rect 2694 2226 2724 2436
rect 2780 2226 2810 2436
rect 2866 2226 2896 2436
rect 2952 2226 2982 2436
rect 3038 2226 3068 2436
rect 3124 2226 3154 2436
rect 3210 2226 3240 2436
rect 3296 2226 3326 2436
rect 3382 2226 3412 2436
rect 3468 2226 3498 2436
rect 3554 2226 3584 2436
rect 4414 2184 4444 2394
rect 4500 2184 4530 2394
rect 5532 2184 5562 2394
rect 5618 2184 5648 2394
rect 6736 2226 6766 2436
rect 6822 2226 6852 2436
rect 7252 2226 7282 2436
rect 7338 2226 7368 2436
rect 7424 2226 7454 2436
rect 7510 2226 7540 2436
rect 7596 2226 7626 2436
rect 7682 2226 7712 2436
rect 7768 2226 7798 2436
rect 7854 2226 7884 2436
rect 7940 2226 7970 2436
rect 8026 2226 8056 2436
rect 8112 2226 8142 2436
rect 8198 2226 8228 2436
rect 8284 2226 8314 2436
rect 8370 2226 8400 2436
rect 8456 2226 8486 2436
rect 8542 2226 8572 2436
rect 8628 2226 8658 2436
rect 8714 2226 8744 2436
rect 8800 2226 8830 2436
rect 8886 2226 8916 2436
rect 8972 2226 9002 2436
rect 9058 2226 9088 2436
rect 9144 2226 9174 2436
rect 9230 2226 9260 2436
rect 9316 2226 9346 2436
rect 9402 2226 9432 2436
rect 9488 2226 9518 2436
rect 9574 2226 9604 2436
rect 9660 2226 9690 2436
rect 9746 2226 9776 2436
rect 9832 2226 9862 2436
rect 9918 2226 9948 2436
rect 10004 2226 10034 2436
rect 10090 2226 10120 2436
rect 10176 2226 10206 2436
rect 10262 2226 10292 2436
rect 10348 2226 10378 2436
rect 10434 2226 10464 2436
rect 10520 2226 10550 2436
rect 10606 2226 10636 2436
rect 10692 2226 10722 2436
rect 10778 2226 10808 2436
rect 10864 2226 10894 2436
rect 10950 2226 10980 2436
rect 11036 2226 11066 2436
rect 11122 2226 11152 2436
rect 11208 2226 11238 2436
rect 11294 2226 11324 2436
rect 200 1791 230 2016
rect 286 1791 316 2016
rect 200 1781 316 1791
rect 200 1747 241 1781
rect 275 1747 316 1781
rect 200 1737 316 1747
rect 372 1791 402 2016
rect 458 1791 488 2016
rect 372 1781 488 1791
rect 372 1747 413 1781
rect 447 1747 488 1781
rect 372 1737 488 1747
rect 544 1791 574 2016
rect 630 1791 660 2016
rect 544 1781 660 1791
rect 544 1747 585 1781
rect 619 1747 660 1781
rect 544 1737 660 1747
rect 716 1791 746 2016
rect 802 1791 832 2016
rect 716 1781 832 1791
rect 716 1747 757 1781
rect 791 1747 832 1781
rect 716 1737 832 1747
rect 888 1791 918 2016
rect 974 1791 1004 2016
rect 888 1781 1004 1791
rect 888 1747 929 1781
rect 963 1747 1004 1781
rect 888 1737 1004 1747
rect 1060 1791 1090 2016
rect 1146 1791 1176 2016
rect 1060 1781 1176 1791
rect 1060 1747 1101 1781
rect 1135 1747 1176 1781
rect 1060 1737 1176 1747
rect 1232 1791 1262 2016
rect 1318 1791 1348 2016
rect 1232 1781 1348 1791
rect 1232 1747 1273 1781
rect 1307 1747 1348 1781
rect 1232 1737 1348 1747
rect 1404 1791 1434 2016
rect 1490 1791 1520 2016
rect 1404 1781 1520 1791
rect 1404 1747 1445 1781
rect 1479 1747 1520 1781
rect 1404 1737 1520 1747
rect 1576 1791 1606 2016
rect 1662 1791 1692 2016
rect 1576 1781 1692 1791
rect 1576 1747 1617 1781
rect 1651 1747 1692 1781
rect 1576 1737 1692 1747
rect 1748 1791 1778 2016
rect 1834 1791 1864 2016
rect 1748 1781 1864 1791
rect 1748 1747 1789 1781
rect 1823 1747 1864 1781
rect 1748 1737 1864 1747
rect 1920 1791 1950 2016
rect 2006 1791 2036 2016
rect 1920 1781 2036 1791
rect 1920 1747 1961 1781
rect 1995 1747 2036 1781
rect 1920 1737 2036 1747
rect 2092 1791 2122 2016
rect 2178 1791 2208 2016
rect 2092 1781 2208 1791
rect 2092 1747 2133 1781
rect 2167 1747 2208 1781
rect 2092 1737 2208 1747
rect 2608 1791 2638 2016
rect 2694 1791 2724 2016
rect 2608 1781 2724 1791
rect 2608 1747 2649 1781
rect 2683 1747 2724 1781
rect 2608 1737 2724 1747
rect 2780 1791 2810 2016
rect 2866 1791 2896 2016
rect 2780 1781 2896 1791
rect 2780 1747 2821 1781
rect 2855 1747 2896 1781
rect 2780 1737 2896 1747
rect 2952 1791 2982 2016
rect 3038 1791 3068 2016
rect 2952 1781 3068 1791
rect 2952 1747 2993 1781
rect 3027 1747 3068 1781
rect 2952 1737 3068 1747
rect 3124 1791 3154 2016
rect 3210 1791 3240 2016
rect 3124 1781 3240 1791
rect 3124 1747 3165 1781
rect 3199 1747 3240 1781
rect 3124 1737 3240 1747
rect 3296 1791 3326 2016
rect 3382 1791 3412 2016
rect 3296 1781 3412 1791
rect 3296 1747 3337 1781
rect 3371 1747 3412 1781
rect 3296 1737 3412 1747
rect 3468 1791 3498 2016
rect 3554 1791 3584 2016
rect 6736 1791 6766 2016
rect 6822 1791 6852 2016
rect 3468 1781 3584 1791
rect 3468 1747 3509 1781
rect 3543 1747 3584 1781
rect 3468 1737 3584 1747
rect 6220 1781 6336 1791
rect 6220 1747 6261 1781
rect 6295 1747 6336 1781
rect 6220 1737 6336 1747
rect 6736 1781 6852 1791
rect 6736 1747 6777 1781
rect 6811 1747 6852 1781
rect 6736 1737 6852 1747
rect 7252 1791 7282 2016
rect 7338 1791 7368 2016
rect 7252 1781 7368 1791
rect 7252 1747 7293 1781
rect 7327 1747 7368 1781
rect 7252 1737 7368 1747
rect 7424 1791 7454 2016
rect 7510 1791 7540 2016
rect 7424 1781 7540 1791
rect 7424 1747 7465 1781
rect 7499 1747 7540 1781
rect 7424 1737 7540 1747
rect 7596 1791 7626 2016
rect 7682 1791 7712 2016
rect 7596 1781 7712 1791
rect 7596 1747 7637 1781
rect 7671 1747 7712 1781
rect 7596 1737 7712 1747
rect 7768 1791 7798 2016
rect 7854 1791 7884 2016
rect 7768 1781 7884 1791
rect 7768 1747 7809 1781
rect 7843 1747 7884 1781
rect 7768 1737 7884 1747
rect 7940 1791 7970 2016
rect 8026 1791 8056 2016
rect 7940 1781 8056 1791
rect 7940 1747 7981 1781
rect 8015 1747 8056 1781
rect 7940 1737 8056 1747
rect 8112 1791 8142 2016
rect 8198 1791 8228 2016
rect 8112 1781 8228 1791
rect 8112 1747 8153 1781
rect 8187 1747 8228 1781
rect 8112 1737 8228 1747
rect 8284 1791 8314 2016
rect 8370 1791 8400 2016
rect 8284 1781 8400 1791
rect 8284 1747 8325 1781
rect 8359 1747 8400 1781
rect 8284 1737 8400 1747
rect 8456 1791 8486 2016
rect 8542 1791 8572 2016
rect 8456 1781 8572 1791
rect 8456 1747 8497 1781
rect 8531 1747 8572 1781
rect 8456 1737 8572 1747
rect 8628 1791 8658 2016
rect 8714 1791 8744 2016
rect 8628 1781 8744 1791
rect 8628 1747 8669 1781
rect 8703 1747 8744 1781
rect 8628 1737 8744 1747
rect 8800 1791 8830 2016
rect 8886 1791 8916 2016
rect 8800 1781 8916 1791
rect 8800 1747 8841 1781
rect 8875 1747 8916 1781
rect 8800 1737 8916 1747
rect 8972 1791 9002 2016
rect 9058 1791 9088 2016
rect 8972 1781 9088 1791
rect 8972 1747 9013 1781
rect 9047 1747 9088 1781
rect 8972 1737 9088 1747
rect 9144 1791 9174 2016
rect 9230 1791 9260 2016
rect 9144 1781 9260 1791
rect 9144 1747 9185 1781
rect 9219 1747 9260 1781
rect 9144 1737 9260 1747
rect 9316 1791 9346 2016
rect 9402 1791 9432 2016
rect 9316 1781 9432 1791
rect 9316 1747 9357 1781
rect 9391 1747 9432 1781
rect 9316 1737 9432 1747
rect 9488 1791 9518 2016
rect 9574 1791 9604 2016
rect 9488 1781 9604 1791
rect 9488 1747 9529 1781
rect 9563 1747 9604 1781
rect 9488 1737 9604 1747
rect 9660 1791 9690 2016
rect 9746 1791 9776 2016
rect 9660 1781 9776 1791
rect 9660 1747 9701 1781
rect 9735 1747 9776 1781
rect 9660 1737 9776 1747
rect 9832 1791 9862 2016
rect 9918 1791 9948 2016
rect 9832 1781 9948 1791
rect 9832 1747 9873 1781
rect 9907 1747 9948 1781
rect 9832 1737 9948 1747
rect 10004 1791 10034 2016
rect 10090 1791 10120 2016
rect 10004 1781 10120 1791
rect 10004 1747 10045 1781
rect 10079 1747 10120 1781
rect 10004 1737 10120 1747
rect 10176 1791 10206 2016
rect 10262 1791 10292 2016
rect 10176 1781 10292 1791
rect 10176 1747 10217 1781
rect 10251 1747 10292 1781
rect 10176 1737 10292 1747
rect 10348 1791 10378 2016
rect 10434 1791 10464 2016
rect 10348 1781 10464 1791
rect 10348 1747 10389 1781
rect 10423 1747 10464 1781
rect 10348 1737 10464 1747
rect 10520 1791 10550 2016
rect 10606 1791 10636 2016
rect 10520 1781 10636 1791
rect 10520 1747 10561 1781
rect 10595 1747 10636 1781
rect 10520 1737 10636 1747
rect 10692 1791 10722 2016
rect 10778 1791 10808 2016
rect 10692 1781 10808 1791
rect 10692 1747 10733 1781
rect 10767 1747 10808 1781
rect 10692 1737 10808 1747
rect 10864 1791 10894 2016
rect 10950 1791 10980 2016
rect 10864 1781 10980 1791
rect 10864 1747 10905 1781
rect 10939 1747 10980 1781
rect 10864 1737 10980 1747
rect 11036 1791 11066 2016
rect 11122 1791 11152 2016
rect 11036 1781 11152 1791
rect 11036 1747 11077 1781
rect 11111 1747 11152 1781
rect 11036 1737 11152 1747
rect 11208 1791 11238 2016
rect 11294 1791 11324 2016
rect 11208 1781 11324 1791
rect 11208 1747 11249 1781
rect 11283 1747 11324 1781
rect 11208 1737 11324 1747
rect 3984 1470 4014 1680
rect 4070 1470 4100 1680
rect 4156 1470 4186 1680
rect 4242 1470 4272 1680
rect 4328 1470 4358 1680
rect 4414 1470 4444 1680
rect 4500 1470 4530 1680
rect 4586 1470 4616 1680
rect 4672 1470 4702 1680
rect 4758 1470 4788 1680
rect 4844 1470 4874 1680
rect 4930 1470 4960 1680
rect 5360 1470 5390 1680
rect 5446 1470 5476 1680
rect 5532 1470 5562 1680
rect 5618 1470 5648 1680
rect 5704 1470 5734 1680
rect 5790 1470 5820 1680
rect 6220 1512 6250 1737
rect 6306 1512 6336 1737
rect 200 1050 230 1260
rect 286 1050 316 1260
rect 372 1050 402 1260
rect 458 1050 488 1260
rect 544 1050 574 1260
rect 630 1050 660 1260
rect 716 1050 746 1260
rect 802 1050 832 1260
rect 888 1050 918 1260
rect 974 1050 1004 1260
rect 1060 1050 1090 1260
rect 1146 1050 1176 1260
rect 1232 1050 1262 1260
rect 1318 1050 1348 1260
rect 1404 1050 1434 1260
rect 1490 1050 1520 1260
rect 1576 1050 1606 1260
rect 1662 1050 1692 1260
rect 1748 1050 1778 1260
rect 1834 1050 1864 1260
rect 1920 1050 1950 1260
rect 2006 1050 2036 1260
rect 2092 1050 2122 1260
rect 2178 1050 2208 1260
rect 2608 1050 2638 1260
rect 2694 1050 2724 1260
rect 2780 1050 2810 1260
rect 2866 1050 2896 1260
rect 2952 1050 2982 1260
rect 3038 1050 3068 1260
rect 3124 1050 3154 1260
rect 3210 1050 3240 1260
rect 3296 1050 3326 1260
rect 3382 1050 3412 1260
rect 3468 1050 3498 1260
rect 3554 1050 3584 1260
rect 3984 1035 4014 1260
rect 4070 1035 4100 1260
rect 3984 1025 4100 1035
rect 3984 991 4025 1025
rect 4059 991 4100 1025
rect 3984 981 4100 991
rect 4156 1035 4186 1260
rect 4242 1035 4272 1260
rect 4156 1025 4272 1035
rect 4156 991 4197 1025
rect 4231 991 4272 1025
rect 4156 981 4272 991
rect 4328 1035 4358 1260
rect 4414 1035 4444 1260
rect 4328 1025 4444 1035
rect 4328 991 4369 1025
rect 4403 991 4444 1025
rect 4328 981 4444 991
rect 4500 1035 4530 1260
rect 4586 1035 4616 1260
rect 4500 1025 4616 1035
rect 4500 991 4541 1025
rect 4575 991 4616 1025
rect 4500 981 4616 991
rect 4672 1035 4702 1260
rect 4758 1035 4788 1260
rect 4672 1025 4788 1035
rect 4672 991 4713 1025
rect 4747 991 4788 1025
rect 4672 981 4788 991
rect 4844 1035 4874 1260
rect 4930 1035 4960 1260
rect 4844 1025 4960 1035
rect 4844 991 4885 1025
rect 4919 991 4960 1025
rect 4844 981 4960 991
rect 5360 1035 5390 1260
rect 5446 1035 5476 1260
rect 5360 1025 5476 1035
rect 5360 991 5401 1025
rect 5435 991 5476 1025
rect 5360 981 5476 991
rect 5532 1035 5562 1260
rect 5618 1035 5648 1260
rect 5532 1025 5648 1035
rect 5532 991 5573 1025
rect 5607 991 5648 1025
rect 5532 981 5648 991
rect 5704 1035 5734 1260
rect 5790 1035 5820 1260
rect 6220 1092 6250 1302
rect 6306 1092 6336 1302
rect 7252 1050 7282 1260
rect 7338 1050 7368 1260
rect 7424 1050 7454 1260
rect 7510 1050 7540 1260
rect 7596 1050 7626 1260
rect 7682 1050 7712 1260
rect 7768 1050 7798 1260
rect 7854 1050 7884 1260
rect 7940 1050 7970 1260
rect 8026 1050 8056 1260
rect 8112 1050 8142 1260
rect 8198 1050 8228 1260
rect 8284 1050 8314 1260
rect 8370 1050 8400 1260
rect 8456 1050 8486 1260
rect 8542 1050 8572 1260
rect 8628 1050 8658 1260
rect 8714 1050 8744 1260
rect 8800 1050 8830 1260
rect 8886 1050 8916 1260
rect 8972 1050 9002 1260
rect 9058 1050 9088 1260
rect 9144 1050 9174 1260
rect 9230 1050 9260 1260
rect 9316 1050 9346 1260
rect 9402 1050 9432 1260
rect 9488 1050 9518 1260
rect 9574 1050 9604 1260
rect 9660 1050 9690 1260
rect 9746 1050 9776 1260
rect 9832 1050 9862 1260
rect 9918 1050 9948 1260
rect 10004 1050 10034 1260
rect 10090 1050 10120 1260
rect 10176 1050 10206 1260
rect 10262 1050 10292 1260
rect 10348 1050 10378 1260
rect 10434 1050 10464 1260
rect 10520 1050 10550 1260
rect 10606 1050 10636 1260
rect 10692 1050 10722 1260
rect 10778 1050 10808 1260
rect 10864 1050 10894 1260
rect 10950 1050 10980 1260
rect 11036 1050 11066 1260
rect 11122 1050 11152 1260
rect 11208 1050 11238 1260
rect 11294 1050 11324 1260
rect 5704 1025 5820 1035
rect 5704 991 5745 1025
rect 5779 991 5820 1025
rect 5704 981 5820 991
rect 200 615 230 840
rect 286 615 316 840
rect 200 605 316 615
rect 200 571 241 605
rect 275 571 316 605
rect 200 561 316 571
rect 372 615 402 840
rect 458 615 488 840
rect 372 605 488 615
rect 372 571 413 605
rect 447 571 488 605
rect 372 561 488 571
rect 544 615 574 840
rect 630 615 660 840
rect 544 605 660 615
rect 544 571 585 605
rect 619 571 660 605
rect 544 561 660 571
rect 716 615 746 840
rect 802 615 832 840
rect 716 605 832 615
rect 716 571 757 605
rect 791 571 832 605
rect 716 561 832 571
rect 888 615 918 840
rect 974 615 1004 840
rect 888 605 1004 615
rect 888 571 929 605
rect 963 571 1004 605
rect 888 561 1004 571
rect 1060 615 1090 840
rect 1146 615 1176 840
rect 1060 605 1176 615
rect 1060 571 1101 605
rect 1135 571 1176 605
rect 1060 561 1176 571
rect 1232 615 1262 840
rect 1318 615 1348 840
rect 1232 605 1348 615
rect 1232 571 1273 605
rect 1307 571 1348 605
rect 1232 561 1348 571
rect 1404 615 1434 840
rect 1490 615 1520 840
rect 1404 605 1520 615
rect 1404 571 1445 605
rect 1479 571 1520 605
rect 1404 561 1520 571
rect 1576 615 1606 840
rect 1662 615 1692 840
rect 1576 605 1692 615
rect 1576 571 1617 605
rect 1651 571 1692 605
rect 1576 561 1692 571
rect 1748 615 1778 840
rect 1834 615 1864 840
rect 1748 605 1864 615
rect 1748 571 1789 605
rect 1823 571 1864 605
rect 1748 561 1864 571
rect 1920 615 1950 840
rect 2006 615 2036 840
rect 1920 605 2036 615
rect 1920 571 1961 605
rect 1995 571 2036 605
rect 1920 561 2036 571
rect 2092 615 2122 840
rect 2178 615 2208 840
rect 2092 605 2208 615
rect 2092 571 2133 605
rect 2167 571 2208 605
rect 2092 561 2208 571
rect 2608 615 2638 840
rect 2694 615 2724 840
rect 2608 605 2724 615
rect 2608 571 2649 605
rect 2683 571 2724 605
rect 2608 561 2724 571
rect 2780 615 2810 840
rect 2866 615 2896 840
rect 2780 605 2896 615
rect 2780 571 2821 605
rect 2855 571 2896 605
rect 2780 561 2896 571
rect 2952 615 2982 840
rect 3038 615 3068 840
rect 2952 605 3068 615
rect 2952 571 2993 605
rect 3027 571 3068 605
rect 2952 561 3068 571
rect 3124 615 3154 840
rect 3210 615 3240 840
rect 3124 605 3240 615
rect 3124 571 3165 605
rect 3199 571 3240 605
rect 3124 561 3240 571
rect 3296 615 3326 840
rect 3382 615 3412 840
rect 3296 605 3412 615
rect 3296 571 3337 605
rect 3371 571 3412 605
rect 3296 561 3412 571
rect 3468 615 3498 840
rect 3554 615 3584 840
rect 3468 605 3584 615
rect 3468 571 3509 605
rect 3543 571 3584 605
rect 3468 561 3584 571
rect 7252 615 7282 840
rect 7338 615 7368 840
rect 7252 605 7368 615
rect 7252 571 7293 605
rect 7327 571 7368 605
rect 7252 561 7368 571
rect 7424 615 7454 840
rect 7510 615 7540 840
rect 7424 605 7540 615
rect 7424 571 7465 605
rect 7499 571 7540 605
rect 7424 561 7540 571
rect 7596 615 7626 840
rect 7682 615 7712 840
rect 7596 605 7712 615
rect 7596 571 7637 605
rect 7671 571 7712 605
rect 7596 561 7712 571
rect 7768 615 7798 840
rect 7854 615 7884 840
rect 7768 605 7884 615
rect 7768 571 7809 605
rect 7843 571 7884 605
rect 7768 561 7884 571
rect 7940 615 7970 840
rect 8026 615 8056 840
rect 7940 605 8056 615
rect 7940 571 7981 605
rect 8015 571 8056 605
rect 7940 561 8056 571
rect 8112 615 8142 840
rect 8198 615 8228 840
rect 8112 605 8228 615
rect 8112 571 8153 605
rect 8187 571 8228 605
rect 8112 561 8228 571
rect 8284 615 8314 840
rect 8370 615 8400 840
rect 8284 605 8400 615
rect 8284 571 8325 605
rect 8359 571 8400 605
rect 8284 561 8400 571
rect 8456 615 8486 840
rect 8542 615 8572 840
rect 8456 605 8572 615
rect 8456 571 8497 605
rect 8531 571 8572 605
rect 8456 561 8572 571
rect 8628 615 8658 840
rect 8714 615 8744 840
rect 8628 605 8744 615
rect 8628 571 8669 605
rect 8703 571 8744 605
rect 8628 561 8744 571
rect 8800 615 8830 840
rect 8886 615 8916 840
rect 8800 605 8916 615
rect 8800 571 8841 605
rect 8875 571 8916 605
rect 8800 561 8916 571
rect 8972 615 9002 840
rect 9058 615 9088 840
rect 8972 605 9088 615
rect 8972 571 9013 605
rect 9047 571 9088 605
rect 8972 561 9088 571
rect 9144 615 9174 840
rect 9230 615 9260 840
rect 9144 605 9260 615
rect 9144 571 9185 605
rect 9219 571 9260 605
rect 9144 561 9260 571
rect 9316 615 9346 840
rect 9402 615 9432 840
rect 9316 605 9432 615
rect 9316 571 9357 605
rect 9391 571 9432 605
rect 9316 561 9432 571
rect 9488 615 9518 840
rect 9574 615 9604 840
rect 9488 605 9604 615
rect 9488 571 9529 605
rect 9563 571 9604 605
rect 9488 561 9604 571
rect 9660 615 9690 840
rect 9746 615 9776 840
rect 9660 605 9776 615
rect 9660 571 9701 605
rect 9735 571 9776 605
rect 9660 561 9776 571
rect 9832 615 9862 840
rect 9918 615 9948 840
rect 9832 605 9948 615
rect 9832 571 9873 605
rect 9907 571 9948 605
rect 9832 561 9948 571
rect 10004 615 10034 840
rect 10090 615 10120 840
rect 10004 605 10120 615
rect 10004 571 10045 605
rect 10079 571 10120 605
rect 10004 561 10120 571
rect 10176 615 10206 840
rect 10262 615 10292 840
rect 10176 605 10292 615
rect 10176 571 10217 605
rect 10251 571 10292 605
rect 10176 561 10292 571
rect 10348 615 10378 840
rect 10434 615 10464 840
rect 10348 605 10464 615
rect 10348 571 10389 605
rect 10423 571 10464 605
rect 10348 561 10464 571
rect 10520 615 10550 840
rect 10606 615 10636 840
rect 10520 605 10636 615
rect 10520 571 10561 605
rect 10595 571 10636 605
rect 10520 561 10636 571
rect 10692 615 10722 840
rect 10778 615 10808 840
rect 10692 605 10808 615
rect 10692 571 10733 605
rect 10767 571 10808 605
rect 10692 561 10808 571
rect 10864 615 10894 840
rect 10950 615 10980 840
rect 10864 605 10980 615
rect 10864 571 10905 605
rect 10939 571 10980 605
rect 10864 561 10980 571
rect 11036 615 11066 840
rect 11122 615 11152 840
rect 11036 605 11152 615
rect 11036 571 11077 605
rect 11111 571 11152 605
rect 11036 561 11152 571
rect 11208 615 11238 840
rect 11294 615 11324 840
rect 11208 605 11324 615
rect 11208 571 11249 605
rect 11283 571 11324 605
rect 11208 561 11324 571
<< polycont >>
rect 1187 3595 1221 3629
rect 3079 3595 3113 3629
rect 6777 3595 6811 3629
rect 9271 3595 9305 3629
rect 6261 3259 6295 3293
rect 4455 2839 4489 2873
rect 5573 2839 5607 2873
rect 241 1747 275 1781
rect 413 1747 447 1781
rect 585 1747 619 1781
rect 757 1747 791 1781
rect 929 1747 963 1781
rect 1101 1747 1135 1781
rect 1273 1747 1307 1781
rect 1445 1747 1479 1781
rect 1617 1747 1651 1781
rect 1789 1747 1823 1781
rect 1961 1747 1995 1781
rect 2133 1747 2167 1781
rect 2649 1747 2683 1781
rect 2821 1747 2855 1781
rect 2993 1747 3027 1781
rect 3165 1747 3199 1781
rect 3337 1747 3371 1781
rect 3509 1747 3543 1781
rect 6261 1747 6295 1781
rect 6777 1747 6811 1781
rect 7293 1747 7327 1781
rect 7465 1747 7499 1781
rect 7637 1747 7671 1781
rect 7809 1747 7843 1781
rect 7981 1747 8015 1781
rect 8153 1747 8187 1781
rect 8325 1747 8359 1781
rect 8497 1747 8531 1781
rect 8669 1747 8703 1781
rect 8841 1747 8875 1781
rect 9013 1747 9047 1781
rect 9185 1747 9219 1781
rect 9357 1747 9391 1781
rect 9529 1747 9563 1781
rect 9701 1747 9735 1781
rect 9873 1747 9907 1781
rect 10045 1747 10079 1781
rect 10217 1747 10251 1781
rect 10389 1747 10423 1781
rect 10561 1747 10595 1781
rect 10733 1747 10767 1781
rect 10905 1747 10939 1781
rect 11077 1747 11111 1781
rect 11249 1747 11283 1781
rect 4025 991 4059 1025
rect 4197 991 4231 1025
rect 4369 991 4403 1025
rect 4541 991 4575 1025
rect 4713 991 4747 1025
rect 4885 991 4919 1025
rect 5401 991 5435 1025
rect 5573 991 5607 1025
rect 5745 991 5779 1025
rect 241 571 275 605
rect 413 571 447 605
rect 585 571 619 605
rect 757 571 791 605
rect 929 571 963 605
rect 1101 571 1135 605
rect 1273 571 1307 605
rect 1445 571 1479 605
rect 1617 571 1651 605
rect 1789 571 1823 605
rect 1961 571 1995 605
rect 2133 571 2167 605
rect 2649 571 2683 605
rect 2821 571 2855 605
rect 2993 571 3027 605
rect 3165 571 3199 605
rect 3337 571 3371 605
rect 3509 571 3543 605
rect 7293 571 7327 605
rect 7465 571 7499 605
rect 7637 571 7671 605
rect 7809 571 7843 605
rect 7981 571 8015 605
rect 8153 571 8187 605
rect 8325 571 8359 605
rect 8497 571 8531 605
rect 8669 571 8703 605
rect 8841 571 8875 605
rect 9013 571 9047 605
rect 9185 571 9219 605
rect 9357 571 9391 605
rect 9529 571 9563 605
rect 9701 571 9735 605
rect 9873 571 9907 605
rect 10045 571 10079 605
rect 10217 571 10251 605
rect 10389 571 10423 605
rect 10561 571 10595 605
rect 10733 571 10767 605
rect 10905 571 10939 605
rect 11077 571 11111 605
rect 11249 571 11283 605
<< locali >>
rect 1179 4049 1229 4133
rect 1179 4015 1187 4049
rect 1221 4015 1229 4049
rect 1179 3931 1229 4015
rect 3071 4049 3121 4133
rect 3071 4015 3079 4049
rect 3113 4015 3121 4049
rect 3071 3931 3121 4015
rect 6769 4049 6819 4133
rect 6769 4015 6777 4049
rect 6811 4015 6819 4049
rect 6769 3931 6819 4015
rect 9263 4049 9313 4133
rect 9263 4015 9271 4049
rect 9305 4015 9313 4049
rect 9263 3931 9313 4015
rect 6253 3713 6303 3797
rect 1179 3629 1229 3713
rect 1179 3595 1187 3629
rect 1221 3595 1229 3629
rect 1179 3511 1229 3595
rect 3071 3629 3121 3713
rect 3071 3595 3079 3629
rect 3113 3595 3121 3629
rect 6253 3679 6261 3713
rect 6295 3679 6303 3713
rect 6253 3595 6303 3679
rect 6769 3629 6819 3713
rect 6769 3595 6777 3629
rect 6811 3595 6819 3629
rect 3071 3511 3121 3595
rect 6769 3511 6819 3595
rect 9263 3629 9313 3713
rect 9263 3595 9271 3629
rect 9305 3595 9313 3629
rect 9263 3511 9313 3595
rect 1093 3336 1143 3461
rect 1093 3302 1101 3336
rect 1135 3302 1143 3336
rect 1093 3268 1143 3302
rect 1093 3234 1101 3268
rect 1135 3234 1143 3268
rect 1093 3200 1143 3234
rect 1093 3166 1101 3200
rect 1135 3166 1143 3200
rect 1093 2873 1143 3166
rect 1093 2839 1101 2873
rect 1135 2839 1143 2873
rect 1093 2755 1143 2839
rect 1179 3336 1229 3461
rect 1179 3302 1187 3336
rect 1221 3302 1229 3336
rect 1179 3268 1229 3302
rect 1179 3234 1187 3268
rect 1221 3234 1229 3268
rect 1179 3200 1229 3234
rect 1179 3166 1187 3200
rect 1221 3166 1229 3200
rect 1179 2789 1229 3166
rect 1179 2755 1187 2789
rect 1221 2755 1229 2789
rect 1265 3336 1315 3461
rect 1265 3302 1273 3336
rect 1307 3302 1315 3336
rect 1265 3268 1315 3302
rect 1265 3234 1273 3268
rect 1307 3234 1315 3268
rect 1265 3200 1315 3234
rect 1265 3166 1273 3200
rect 1307 3166 1315 3200
rect 1265 2873 1315 3166
rect 1265 2839 1273 2873
rect 1307 2839 1315 2873
rect 1265 2755 1315 2839
rect 2985 3336 3035 3461
rect 2985 3302 2993 3336
rect 3027 3302 3035 3336
rect 2985 3268 3035 3302
rect 2985 3234 2993 3268
rect 3027 3234 3035 3268
rect 2985 3200 3035 3234
rect 2985 3166 2993 3200
rect 3027 3166 3035 3200
rect 2985 2873 3035 3166
rect 2985 2839 2993 2873
rect 3027 2839 3035 2873
rect 2985 2755 3035 2839
rect 3071 3336 3121 3461
rect 3071 3302 3079 3336
rect 3113 3302 3121 3336
rect 3071 3268 3121 3302
rect 3071 3234 3079 3268
rect 3113 3234 3121 3268
rect 3071 3200 3121 3234
rect 3071 3166 3079 3200
rect 3113 3166 3121 3200
rect 3071 2789 3121 3166
rect 3071 2755 3079 2789
rect 3113 2755 3121 2789
rect 3157 3336 3207 3461
rect 3157 3302 3165 3336
rect 3199 3302 3207 3336
rect 3157 3268 3207 3302
rect 3157 3234 3165 3268
rect 3199 3234 3207 3268
rect 3157 3200 3207 3234
rect 3157 3166 3165 3200
rect 3199 3166 3207 3200
rect 4447 3293 4497 3377
rect 4447 3259 4455 3293
rect 4489 3259 4497 3293
rect 4447 3175 4497 3259
rect 5565 3293 5615 3377
rect 5565 3259 5573 3293
rect 5607 3259 5615 3293
rect 5565 3175 5615 3259
rect 6253 3293 6303 3377
rect 6683 3336 6733 3461
rect 6683 3302 6691 3336
rect 6725 3302 6733 3336
rect 6253 3259 6261 3293
rect 6295 3259 6303 3293
rect 6253 3175 6303 3259
rect 6597 3259 6605 3293
rect 6639 3259 6647 3293
rect 3157 2873 3207 3166
rect 6167 3000 6217 3125
rect 6167 2966 6175 3000
rect 6209 2966 6217 3000
rect 3157 2839 3165 2873
rect 3199 2839 3207 2873
rect 3157 2755 3207 2839
rect 4447 2873 4497 2957
rect 4447 2839 4455 2873
rect 4489 2839 4497 2873
rect 4447 2755 4497 2839
rect 5565 2873 5615 2957
rect 5565 2839 5573 2873
rect 5607 2839 5615 2873
rect 5565 2755 5615 2839
rect 6167 2932 6217 2966
rect 6167 2898 6175 2932
rect 6209 2898 6217 2932
rect 6167 2864 6217 2898
rect 6167 2830 6175 2864
rect 6209 2830 6217 2864
rect 147 2537 197 2621
rect 147 2503 155 2537
rect 189 2503 197 2537
rect 147 2210 197 2503
rect 147 2176 155 2210
rect 189 2176 197 2210
rect 147 2142 197 2176
rect 147 2108 155 2142
rect 189 2108 197 2142
rect 147 2074 197 2108
rect 147 2040 155 2074
rect 189 2040 197 2074
rect 147 1915 197 2040
rect 233 2587 241 2621
rect 275 2587 283 2621
rect 233 2210 283 2587
rect 233 2176 241 2210
rect 275 2176 283 2210
rect 233 2142 283 2176
rect 233 2108 241 2142
rect 275 2108 283 2142
rect 233 2074 283 2108
rect 233 2040 241 2074
rect 275 2040 283 2074
rect 233 1915 283 2040
rect 319 2537 369 2621
rect 319 2503 327 2537
rect 361 2503 369 2537
rect 319 2210 369 2503
rect 319 2176 327 2210
rect 361 2176 369 2210
rect 319 2142 369 2176
rect 319 2108 327 2142
rect 361 2108 369 2142
rect 319 2074 369 2108
rect 319 2040 327 2074
rect 361 2040 369 2074
rect 319 1915 369 2040
rect 405 2587 413 2621
rect 447 2587 455 2621
rect 405 2210 455 2587
rect 405 2176 413 2210
rect 447 2176 455 2210
rect 405 2142 455 2176
rect 405 2108 413 2142
rect 447 2108 455 2142
rect 405 2074 455 2108
rect 405 2040 413 2074
rect 447 2040 455 2074
rect 405 1915 455 2040
rect 491 2537 541 2621
rect 491 2503 499 2537
rect 533 2503 541 2537
rect 491 2210 541 2503
rect 491 2176 499 2210
rect 533 2176 541 2210
rect 491 2142 541 2176
rect 491 2108 499 2142
rect 533 2108 541 2142
rect 491 2074 541 2108
rect 491 2040 499 2074
rect 533 2040 541 2074
rect 491 1915 541 2040
rect 577 2587 585 2621
rect 619 2587 627 2621
rect 577 2210 627 2587
rect 577 2176 585 2210
rect 619 2176 627 2210
rect 577 2142 627 2176
rect 577 2108 585 2142
rect 619 2108 627 2142
rect 577 2074 627 2108
rect 577 2040 585 2074
rect 619 2040 627 2074
rect 577 1915 627 2040
rect 663 2537 713 2621
rect 663 2503 671 2537
rect 705 2503 713 2537
rect 663 2210 713 2503
rect 663 2176 671 2210
rect 705 2176 713 2210
rect 663 2142 713 2176
rect 663 2108 671 2142
rect 705 2108 713 2142
rect 663 2074 713 2108
rect 663 2040 671 2074
rect 705 2040 713 2074
rect 663 1915 713 2040
rect 749 2587 757 2621
rect 791 2587 799 2621
rect 749 2210 799 2587
rect 749 2176 757 2210
rect 791 2176 799 2210
rect 749 2142 799 2176
rect 749 2108 757 2142
rect 791 2108 799 2142
rect 749 2074 799 2108
rect 749 2040 757 2074
rect 791 2040 799 2074
rect 749 1915 799 2040
rect 835 2537 885 2621
rect 835 2503 843 2537
rect 877 2503 885 2537
rect 835 2210 885 2503
rect 835 2176 843 2210
rect 877 2176 885 2210
rect 835 2142 885 2176
rect 835 2108 843 2142
rect 877 2108 885 2142
rect 835 2074 885 2108
rect 835 2040 843 2074
rect 877 2040 885 2074
rect 835 1915 885 2040
rect 921 2587 929 2621
rect 963 2587 971 2621
rect 921 2210 971 2587
rect 921 2176 929 2210
rect 963 2176 971 2210
rect 921 2142 971 2176
rect 921 2108 929 2142
rect 963 2108 971 2142
rect 921 2074 971 2108
rect 921 2040 929 2074
rect 963 2040 971 2074
rect 921 1915 971 2040
rect 1007 2537 1057 2621
rect 1007 2503 1015 2537
rect 1049 2503 1057 2537
rect 1007 2210 1057 2503
rect 1007 2176 1015 2210
rect 1049 2176 1057 2210
rect 1007 2142 1057 2176
rect 1007 2108 1015 2142
rect 1049 2108 1057 2142
rect 1007 2074 1057 2108
rect 1007 2040 1015 2074
rect 1049 2040 1057 2074
rect 1007 1915 1057 2040
rect 1093 2587 1101 2621
rect 1135 2587 1143 2621
rect 1093 2210 1143 2587
rect 1093 2176 1101 2210
rect 1135 2176 1143 2210
rect 1093 2142 1143 2176
rect 1093 2108 1101 2142
rect 1135 2108 1143 2142
rect 1093 2074 1143 2108
rect 1093 2040 1101 2074
rect 1135 2040 1143 2074
rect 1093 1915 1143 2040
rect 1179 2537 1229 2621
rect 1179 2503 1187 2537
rect 1221 2503 1229 2537
rect 1179 2210 1229 2503
rect 1179 2176 1187 2210
rect 1221 2176 1229 2210
rect 1179 2142 1229 2176
rect 1179 2108 1187 2142
rect 1221 2108 1229 2142
rect 1179 2074 1229 2108
rect 1179 2040 1187 2074
rect 1221 2040 1229 2074
rect 1179 1915 1229 2040
rect 1265 2587 1273 2621
rect 1307 2587 1315 2621
rect 1265 2210 1315 2587
rect 1265 2176 1273 2210
rect 1307 2176 1315 2210
rect 1265 2142 1315 2176
rect 1265 2108 1273 2142
rect 1307 2108 1315 2142
rect 1265 2074 1315 2108
rect 1265 2040 1273 2074
rect 1307 2040 1315 2074
rect 1265 1915 1315 2040
rect 1351 2537 1401 2621
rect 1351 2503 1359 2537
rect 1393 2503 1401 2537
rect 1351 2210 1401 2503
rect 1351 2176 1359 2210
rect 1393 2176 1401 2210
rect 1351 2142 1401 2176
rect 1351 2108 1359 2142
rect 1393 2108 1401 2142
rect 1351 2074 1401 2108
rect 1351 2040 1359 2074
rect 1393 2040 1401 2074
rect 1351 1915 1401 2040
rect 1437 2587 1445 2621
rect 1479 2587 1487 2621
rect 1437 2210 1487 2587
rect 1437 2176 1445 2210
rect 1479 2176 1487 2210
rect 1437 2142 1487 2176
rect 1437 2108 1445 2142
rect 1479 2108 1487 2142
rect 1437 2074 1487 2108
rect 1437 2040 1445 2074
rect 1479 2040 1487 2074
rect 1437 1915 1487 2040
rect 1523 2537 1573 2621
rect 1523 2503 1531 2537
rect 1565 2503 1573 2537
rect 1523 2210 1573 2503
rect 1523 2176 1531 2210
rect 1565 2176 1573 2210
rect 1523 2142 1573 2176
rect 1523 2108 1531 2142
rect 1565 2108 1573 2142
rect 1523 2074 1573 2108
rect 1523 2040 1531 2074
rect 1565 2040 1573 2074
rect 1523 1915 1573 2040
rect 1609 2587 1617 2621
rect 1651 2587 1659 2621
rect 1609 2210 1659 2587
rect 1609 2176 1617 2210
rect 1651 2176 1659 2210
rect 1609 2142 1659 2176
rect 1609 2108 1617 2142
rect 1651 2108 1659 2142
rect 1609 2074 1659 2108
rect 1609 2040 1617 2074
rect 1651 2040 1659 2074
rect 1609 1915 1659 2040
rect 1695 2537 1745 2621
rect 1695 2503 1703 2537
rect 1737 2503 1745 2537
rect 1695 2210 1745 2503
rect 1695 2176 1703 2210
rect 1737 2176 1745 2210
rect 1695 2142 1745 2176
rect 1695 2108 1703 2142
rect 1737 2108 1745 2142
rect 1695 2074 1745 2108
rect 1695 2040 1703 2074
rect 1737 2040 1745 2074
rect 1695 1915 1745 2040
rect 1781 2587 1789 2621
rect 1823 2587 1831 2621
rect 1781 2210 1831 2587
rect 1781 2176 1789 2210
rect 1823 2176 1831 2210
rect 1781 2142 1831 2176
rect 1781 2108 1789 2142
rect 1823 2108 1831 2142
rect 1781 2074 1831 2108
rect 1781 2040 1789 2074
rect 1823 2040 1831 2074
rect 1781 1915 1831 2040
rect 1867 2537 1917 2621
rect 1867 2503 1875 2537
rect 1909 2503 1917 2537
rect 1867 2210 1917 2503
rect 1867 2176 1875 2210
rect 1909 2176 1917 2210
rect 1867 2142 1917 2176
rect 1867 2108 1875 2142
rect 1909 2108 1917 2142
rect 1867 2074 1917 2108
rect 1867 2040 1875 2074
rect 1909 2040 1917 2074
rect 1867 1915 1917 2040
rect 1953 2587 1961 2621
rect 1995 2587 2003 2621
rect 1953 2210 2003 2587
rect 1953 2176 1961 2210
rect 1995 2176 2003 2210
rect 1953 2142 2003 2176
rect 1953 2108 1961 2142
rect 1995 2108 2003 2142
rect 1953 2074 2003 2108
rect 1953 2040 1961 2074
rect 1995 2040 2003 2074
rect 1953 1915 2003 2040
rect 2039 2537 2089 2621
rect 2039 2503 2047 2537
rect 2081 2503 2089 2537
rect 2039 2210 2089 2503
rect 2039 2176 2047 2210
rect 2081 2176 2089 2210
rect 2039 2142 2089 2176
rect 2039 2108 2047 2142
rect 2081 2108 2089 2142
rect 2039 2074 2089 2108
rect 2039 2040 2047 2074
rect 2081 2040 2089 2074
rect 2039 1915 2089 2040
rect 2125 2587 2133 2621
rect 2167 2587 2175 2621
rect 2125 2210 2175 2587
rect 2125 2176 2133 2210
rect 2167 2176 2175 2210
rect 2125 2142 2175 2176
rect 2125 2108 2133 2142
rect 2167 2108 2175 2142
rect 2125 2074 2175 2108
rect 2125 2040 2133 2074
rect 2167 2040 2175 2074
rect 2125 1915 2175 2040
rect 2211 2537 2261 2621
rect 2211 2503 2219 2537
rect 2253 2503 2261 2537
rect 2211 2210 2261 2503
rect 2211 2176 2219 2210
rect 2253 2176 2261 2210
rect 2211 2142 2261 2176
rect 2211 2108 2219 2142
rect 2253 2108 2261 2142
rect 2211 2074 2261 2108
rect 2211 2040 2219 2074
rect 2253 2040 2261 2074
rect 2211 1915 2261 2040
rect 2555 2537 2605 2621
rect 2555 2503 2563 2537
rect 2597 2503 2605 2537
rect 2555 2210 2605 2503
rect 2555 2176 2563 2210
rect 2597 2176 2605 2210
rect 2555 2142 2605 2176
rect 2555 2108 2563 2142
rect 2597 2108 2605 2142
rect 2555 2074 2605 2108
rect 2555 2040 2563 2074
rect 2597 2040 2605 2074
rect 2555 1915 2605 2040
rect 2641 2587 2649 2621
rect 2683 2587 2691 2621
rect 2641 2210 2691 2587
rect 2641 2176 2649 2210
rect 2683 2176 2691 2210
rect 2641 2142 2691 2176
rect 2641 2108 2649 2142
rect 2683 2108 2691 2142
rect 2641 2074 2691 2108
rect 2641 2040 2649 2074
rect 2683 2040 2691 2074
rect 2641 1915 2691 2040
rect 2727 2537 2777 2621
rect 2727 2503 2735 2537
rect 2769 2503 2777 2537
rect 2727 2210 2777 2503
rect 2727 2176 2735 2210
rect 2769 2176 2777 2210
rect 2727 2142 2777 2176
rect 2727 2108 2735 2142
rect 2769 2108 2777 2142
rect 2727 2074 2777 2108
rect 2727 2040 2735 2074
rect 2769 2040 2777 2074
rect 2727 1915 2777 2040
rect 2813 2587 2821 2621
rect 2855 2587 2863 2621
rect 2813 2210 2863 2587
rect 2813 2176 2821 2210
rect 2855 2176 2863 2210
rect 2813 2142 2863 2176
rect 2813 2108 2821 2142
rect 2855 2108 2863 2142
rect 2813 2074 2863 2108
rect 2813 2040 2821 2074
rect 2855 2040 2863 2074
rect 2813 1915 2863 2040
rect 2899 2537 2949 2621
rect 2899 2503 2907 2537
rect 2941 2503 2949 2537
rect 2899 2210 2949 2503
rect 2899 2176 2907 2210
rect 2941 2176 2949 2210
rect 2899 2142 2949 2176
rect 2899 2108 2907 2142
rect 2941 2108 2949 2142
rect 2899 2074 2949 2108
rect 2899 2040 2907 2074
rect 2941 2040 2949 2074
rect 2899 1915 2949 2040
rect 2985 2587 2993 2621
rect 3027 2587 3035 2621
rect 2985 2210 3035 2587
rect 2985 2176 2993 2210
rect 3027 2176 3035 2210
rect 2985 2142 3035 2176
rect 2985 2108 2993 2142
rect 3027 2108 3035 2142
rect 2985 2074 3035 2108
rect 2985 2040 2993 2074
rect 3027 2040 3035 2074
rect 2985 1915 3035 2040
rect 3071 2537 3121 2621
rect 3071 2503 3079 2537
rect 3113 2503 3121 2537
rect 3071 2210 3121 2503
rect 3071 2176 3079 2210
rect 3113 2176 3121 2210
rect 3071 2142 3121 2176
rect 3071 2108 3079 2142
rect 3113 2108 3121 2142
rect 3071 2074 3121 2108
rect 3071 2040 3079 2074
rect 3113 2040 3121 2074
rect 3071 1915 3121 2040
rect 3157 2587 3165 2621
rect 3199 2587 3207 2621
rect 3157 2210 3207 2587
rect 3157 2176 3165 2210
rect 3199 2176 3207 2210
rect 3157 2142 3207 2176
rect 3157 2108 3165 2142
rect 3199 2108 3207 2142
rect 3157 2074 3207 2108
rect 3157 2040 3165 2074
rect 3199 2040 3207 2074
rect 3157 1915 3207 2040
rect 3243 2537 3293 2621
rect 3243 2503 3251 2537
rect 3285 2503 3293 2537
rect 3243 2210 3293 2503
rect 3243 2176 3251 2210
rect 3285 2176 3293 2210
rect 3243 2142 3293 2176
rect 3243 2108 3251 2142
rect 3285 2108 3293 2142
rect 3243 2074 3293 2108
rect 3243 2040 3251 2074
rect 3285 2040 3293 2074
rect 3243 1915 3293 2040
rect 3329 2587 3337 2621
rect 3371 2587 3379 2621
rect 3329 2210 3379 2587
rect 3329 2176 3337 2210
rect 3371 2176 3379 2210
rect 3329 2142 3379 2176
rect 3329 2108 3337 2142
rect 3371 2108 3379 2142
rect 3329 2074 3379 2108
rect 3329 2040 3337 2074
rect 3371 2040 3379 2074
rect 3329 1915 3379 2040
rect 3415 2537 3465 2621
rect 3415 2503 3423 2537
rect 3457 2503 3465 2537
rect 3415 2210 3465 2503
rect 3415 2176 3423 2210
rect 3457 2176 3465 2210
rect 3415 2142 3465 2176
rect 3415 2108 3423 2142
rect 3457 2108 3465 2142
rect 3415 2074 3465 2108
rect 3415 2040 3423 2074
rect 3457 2040 3465 2074
rect 3415 1915 3465 2040
rect 3501 2587 3509 2621
rect 3543 2587 3551 2621
rect 3501 2210 3551 2587
rect 3501 2176 3509 2210
rect 3543 2176 3551 2210
rect 3501 2142 3551 2176
rect 3501 2108 3509 2142
rect 3543 2108 3551 2142
rect 3501 2074 3551 2108
rect 3501 2040 3509 2074
rect 3543 2040 3551 2074
rect 3501 1915 3551 2040
rect 3587 2537 3637 2621
rect 3587 2503 3595 2537
rect 3629 2503 3637 2537
rect 3587 2210 3637 2503
rect 3587 2176 3595 2210
rect 3629 2176 3637 2210
rect 3587 2142 3637 2176
rect 3587 2108 3595 2142
rect 3629 2108 3637 2142
rect 3587 2074 3637 2108
rect 3587 2040 3595 2074
rect 3629 2040 3637 2074
rect 3587 1915 3637 2040
rect 4361 2580 4411 2705
rect 4361 2546 4369 2580
rect 4403 2546 4411 2580
rect 4361 2512 4411 2546
rect 4361 2478 4369 2512
rect 4403 2478 4411 2512
rect 4361 2444 4411 2478
rect 4361 2410 4369 2444
rect 4403 2410 4411 2444
rect 4361 2117 4411 2410
rect 4361 2083 4369 2117
rect 4403 2083 4411 2117
rect 4361 1999 4411 2083
rect 4447 2580 4497 2705
rect 4447 2546 4455 2580
rect 4489 2546 4497 2580
rect 4447 2512 4497 2546
rect 4447 2478 4455 2512
rect 4489 2478 4497 2512
rect 4447 2444 4497 2478
rect 4447 2410 4455 2444
rect 4489 2410 4497 2444
rect 4447 2033 4497 2410
rect 4447 1999 4455 2033
rect 4489 1999 4497 2033
rect 4533 2580 4583 2705
rect 4533 2546 4541 2580
rect 4575 2546 4583 2580
rect 4533 2512 4583 2546
rect 4533 2478 4541 2512
rect 4575 2478 4583 2512
rect 4533 2444 4583 2478
rect 4533 2410 4541 2444
rect 4575 2410 4583 2444
rect 4533 2117 4583 2410
rect 4533 2083 4541 2117
rect 4575 2083 4583 2117
rect 4533 1999 4583 2083
rect 5479 2580 5529 2705
rect 5479 2546 5487 2580
rect 5521 2546 5529 2580
rect 5479 2512 5529 2546
rect 5479 2478 5487 2512
rect 5521 2478 5529 2512
rect 5479 2444 5529 2478
rect 5479 2410 5487 2444
rect 5521 2410 5529 2444
rect 5479 2117 5529 2410
rect 5479 2083 5487 2117
rect 5521 2083 5529 2117
rect 5479 1999 5529 2083
rect 5565 2580 5615 2705
rect 5565 2546 5573 2580
rect 5607 2546 5615 2580
rect 5565 2512 5615 2546
rect 5565 2478 5573 2512
rect 5607 2478 5615 2512
rect 5565 2444 5615 2478
rect 5565 2410 5573 2444
rect 5607 2410 5615 2444
rect 5565 2033 5615 2410
rect 5565 1999 5573 2033
rect 5607 1999 5615 2033
rect 5651 2580 5701 2705
rect 5651 2546 5659 2580
rect 5693 2546 5701 2580
rect 5651 2512 5701 2546
rect 5651 2478 5659 2512
rect 5693 2478 5701 2512
rect 5651 2444 5701 2478
rect 5651 2410 5659 2444
rect 5693 2410 5701 2444
rect 6167 2537 6217 2830
rect 6167 2503 6175 2537
rect 6209 2503 6217 2537
rect 6167 2419 6217 2503
rect 6253 3000 6303 3125
rect 6253 2966 6261 3000
rect 6295 2966 6303 3000
rect 6253 2932 6303 2966
rect 6253 2898 6261 2932
rect 6295 2898 6303 2932
rect 6253 2864 6303 2898
rect 6253 2830 6261 2864
rect 6295 2830 6303 2864
rect 6253 2453 6303 2830
rect 6253 2419 6261 2453
rect 6295 2419 6303 2453
rect 6339 3000 6389 3125
rect 6339 2966 6347 3000
rect 6381 2966 6389 3000
rect 6339 2932 6389 2966
rect 6339 2898 6347 2932
rect 6381 2898 6389 2932
rect 6339 2864 6389 2898
rect 6339 2830 6347 2864
rect 6381 2830 6389 2864
rect 6339 2537 6389 2830
rect 6597 2789 6647 3259
rect 6597 2755 6605 2789
rect 6639 2755 6647 2789
rect 6683 3268 6733 3302
rect 6683 3234 6691 3268
rect 6725 3234 6733 3268
rect 6683 3200 6733 3234
rect 6683 3166 6691 3200
rect 6725 3166 6733 3200
rect 6683 2873 6733 3166
rect 6683 2839 6691 2873
rect 6725 2839 6733 2873
rect 6683 2755 6733 2839
rect 6769 3336 6819 3461
rect 6769 3302 6777 3336
rect 6811 3302 6819 3336
rect 6769 3268 6819 3302
rect 6769 3234 6777 3268
rect 6811 3234 6819 3268
rect 6769 3200 6819 3234
rect 6769 3166 6777 3200
rect 6811 3166 6819 3200
rect 6769 2789 6819 3166
rect 6769 2755 6777 2789
rect 6811 2755 6819 2789
rect 6855 3336 6905 3461
rect 6855 3302 6863 3336
rect 6897 3302 6905 3336
rect 6855 3268 6905 3302
rect 6855 3234 6863 3268
rect 6897 3234 6905 3268
rect 6855 3200 6905 3234
rect 6855 3166 6863 3200
rect 6897 3166 6905 3200
rect 6855 2873 6905 3166
rect 6855 2839 6863 2873
rect 6897 2839 6905 2873
rect 6855 2755 6905 2839
rect 9177 3336 9227 3461
rect 9177 3302 9185 3336
rect 9219 3302 9227 3336
rect 9177 3268 9227 3302
rect 9177 3234 9185 3268
rect 9219 3234 9227 3268
rect 9177 3200 9227 3234
rect 9177 3166 9185 3200
rect 9219 3166 9227 3200
rect 9177 2873 9227 3166
rect 9177 2839 9185 2873
rect 9219 2839 9227 2873
rect 9177 2755 9227 2839
rect 9263 3336 9313 3461
rect 9263 3302 9271 3336
rect 9305 3302 9313 3336
rect 9263 3268 9313 3302
rect 9263 3234 9271 3268
rect 9305 3234 9313 3268
rect 9263 3200 9313 3234
rect 9263 3166 9271 3200
rect 9305 3166 9313 3200
rect 9263 2789 9313 3166
rect 9263 2755 9271 2789
rect 9305 2755 9313 2789
rect 9349 3336 9399 3461
rect 9349 3302 9357 3336
rect 9391 3302 9399 3336
rect 9349 3268 9399 3302
rect 9349 3234 9357 3268
rect 9391 3234 9399 3268
rect 9349 3200 9399 3234
rect 9349 3166 9357 3200
rect 9391 3166 9399 3200
rect 9349 2873 9399 3166
rect 9349 2839 9357 2873
rect 9391 2839 9399 2873
rect 9349 2755 9399 2839
rect 6597 2621 6647 2755
rect 6597 2587 6605 2621
rect 6639 2587 6647 2621
rect 6339 2503 6347 2537
rect 6381 2503 6389 2537
rect 6339 2419 6389 2503
rect 6683 2537 6733 2621
rect 6683 2503 6691 2537
rect 6725 2503 6733 2537
rect 5651 2117 5701 2410
rect 5651 2083 5659 2117
rect 5693 2083 5701 2117
rect 6253 2201 6303 2285
rect 6253 2167 6261 2201
rect 6295 2167 6303 2201
rect 6253 2083 6303 2167
rect 6683 2210 6733 2503
rect 6683 2176 6691 2210
rect 6725 2176 6733 2210
rect 6683 2142 6733 2176
rect 6683 2108 6691 2142
rect 6725 2108 6733 2142
rect 5651 1999 5701 2083
rect 6683 2074 6733 2108
rect 6683 2040 6691 2074
rect 6725 2040 6733 2074
rect 5221 1915 5229 1949
rect 5263 1915 5271 1949
rect 6683 1915 6733 2040
rect 6769 2587 6777 2621
rect 6811 2587 6819 2621
rect 6769 2210 6819 2587
rect 6769 2176 6777 2210
rect 6811 2176 6819 2210
rect 6769 2142 6819 2176
rect 6769 2108 6777 2142
rect 6811 2108 6819 2142
rect 6769 2074 6819 2108
rect 6769 2040 6777 2074
rect 6811 2040 6819 2074
rect 6769 1915 6819 2040
rect 6855 2537 6905 2621
rect 6855 2503 6863 2537
rect 6897 2503 6905 2537
rect 6855 2210 6905 2503
rect 6855 2176 6863 2210
rect 6897 2176 6905 2210
rect 6855 2142 6905 2176
rect 6855 2108 6863 2142
rect 6897 2108 6905 2142
rect 6855 2074 6905 2108
rect 6855 2040 6863 2074
rect 6897 2040 6905 2074
rect 6855 1915 6905 2040
rect 7199 2537 7249 2621
rect 7199 2503 7207 2537
rect 7241 2503 7249 2537
rect 7199 2210 7249 2503
rect 7199 2176 7207 2210
rect 7241 2176 7249 2210
rect 7199 2142 7249 2176
rect 7199 2108 7207 2142
rect 7241 2108 7249 2142
rect 7199 2074 7249 2108
rect 7199 2040 7207 2074
rect 7241 2040 7249 2074
rect 7199 1915 7249 2040
rect 7285 2587 7293 2621
rect 7327 2587 7335 2621
rect 7285 2210 7335 2587
rect 7285 2176 7293 2210
rect 7327 2176 7335 2210
rect 7285 2142 7335 2176
rect 7285 2108 7293 2142
rect 7327 2108 7335 2142
rect 7285 2074 7335 2108
rect 7285 2040 7293 2074
rect 7327 2040 7335 2074
rect 7285 1915 7335 2040
rect 7371 2537 7421 2621
rect 7371 2503 7379 2537
rect 7413 2503 7421 2537
rect 7371 2210 7421 2503
rect 7371 2176 7379 2210
rect 7413 2176 7421 2210
rect 7371 2142 7421 2176
rect 7371 2108 7379 2142
rect 7413 2108 7421 2142
rect 7371 2074 7421 2108
rect 7371 2040 7379 2074
rect 7413 2040 7421 2074
rect 7371 1915 7421 2040
rect 7457 2587 7465 2621
rect 7499 2587 7507 2621
rect 7457 2210 7507 2587
rect 7457 2176 7465 2210
rect 7499 2176 7507 2210
rect 7457 2142 7507 2176
rect 7457 2108 7465 2142
rect 7499 2108 7507 2142
rect 7457 2074 7507 2108
rect 7457 2040 7465 2074
rect 7499 2040 7507 2074
rect 7457 1915 7507 2040
rect 7543 2537 7593 2621
rect 7543 2503 7551 2537
rect 7585 2503 7593 2537
rect 7543 2210 7593 2503
rect 7543 2176 7551 2210
rect 7585 2176 7593 2210
rect 7543 2142 7593 2176
rect 7543 2108 7551 2142
rect 7585 2108 7593 2142
rect 7543 2074 7593 2108
rect 7543 2040 7551 2074
rect 7585 2040 7593 2074
rect 7543 1915 7593 2040
rect 7629 2587 7637 2621
rect 7671 2587 7679 2621
rect 7629 2210 7679 2587
rect 7629 2176 7637 2210
rect 7671 2176 7679 2210
rect 7629 2142 7679 2176
rect 7629 2108 7637 2142
rect 7671 2108 7679 2142
rect 7629 2074 7679 2108
rect 7629 2040 7637 2074
rect 7671 2040 7679 2074
rect 7629 1915 7679 2040
rect 7715 2537 7765 2621
rect 7715 2503 7723 2537
rect 7757 2503 7765 2537
rect 7715 2210 7765 2503
rect 7715 2176 7723 2210
rect 7757 2176 7765 2210
rect 7715 2142 7765 2176
rect 7715 2108 7723 2142
rect 7757 2108 7765 2142
rect 7715 2074 7765 2108
rect 7715 2040 7723 2074
rect 7757 2040 7765 2074
rect 7715 1915 7765 2040
rect 7801 2587 7809 2621
rect 7843 2587 7851 2621
rect 7801 2210 7851 2587
rect 7801 2176 7809 2210
rect 7843 2176 7851 2210
rect 7801 2142 7851 2176
rect 7801 2108 7809 2142
rect 7843 2108 7851 2142
rect 7801 2074 7851 2108
rect 7801 2040 7809 2074
rect 7843 2040 7851 2074
rect 7801 1915 7851 2040
rect 7887 2537 7937 2621
rect 7887 2503 7895 2537
rect 7929 2503 7937 2537
rect 7887 2210 7937 2503
rect 7887 2176 7895 2210
rect 7929 2176 7937 2210
rect 7887 2142 7937 2176
rect 7887 2108 7895 2142
rect 7929 2108 7937 2142
rect 7887 2074 7937 2108
rect 7887 2040 7895 2074
rect 7929 2040 7937 2074
rect 7887 1915 7937 2040
rect 7973 2587 7981 2621
rect 8015 2587 8023 2621
rect 7973 2210 8023 2587
rect 7973 2176 7981 2210
rect 8015 2176 8023 2210
rect 7973 2142 8023 2176
rect 7973 2108 7981 2142
rect 8015 2108 8023 2142
rect 7973 2074 8023 2108
rect 7973 2040 7981 2074
rect 8015 2040 8023 2074
rect 7973 1915 8023 2040
rect 8059 2537 8109 2621
rect 8059 2503 8067 2537
rect 8101 2503 8109 2537
rect 8059 2210 8109 2503
rect 8059 2176 8067 2210
rect 8101 2176 8109 2210
rect 8059 2142 8109 2176
rect 8059 2108 8067 2142
rect 8101 2108 8109 2142
rect 8059 2074 8109 2108
rect 8059 2040 8067 2074
rect 8101 2040 8109 2074
rect 8059 1915 8109 2040
rect 8145 2587 8153 2621
rect 8187 2587 8195 2621
rect 8145 2210 8195 2587
rect 8145 2176 8153 2210
rect 8187 2176 8195 2210
rect 8145 2142 8195 2176
rect 8145 2108 8153 2142
rect 8187 2108 8195 2142
rect 8145 2074 8195 2108
rect 8145 2040 8153 2074
rect 8187 2040 8195 2074
rect 8145 1915 8195 2040
rect 8231 2537 8281 2621
rect 8231 2503 8239 2537
rect 8273 2503 8281 2537
rect 8231 2210 8281 2503
rect 8231 2176 8239 2210
rect 8273 2176 8281 2210
rect 8231 2142 8281 2176
rect 8231 2108 8239 2142
rect 8273 2108 8281 2142
rect 8231 2074 8281 2108
rect 8231 2040 8239 2074
rect 8273 2040 8281 2074
rect 8231 1915 8281 2040
rect 8317 2587 8325 2621
rect 8359 2587 8367 2621
rect 8317 2210 8367 2587
rect 8317 2176 8325 2210
rect 8359 2176 8367 2210
rect 8317 2142 8367 2176
rect 8317 2108 8325 2142
rect 8359 2108 8367 2142
rect 8317 2074 8367 2108
rect 8317 2040 8325 2074
rect 8359 2040 8367 2074
rect 8317 1915 8367 2040
rect 8403 2537 8453 2621
rect 8403 2503 8411 2537
rect 8445 2503 8453 2537
rect 8403 2210 8453 2503
rect 8403 2176 8411 2210
rect 8445 2176 8453 2210
rect 8403 2142 8453 2176
rect 8403 2108 8411 2142
rect 8445 2108 8453 2142
rect 8403 2074 8453 2108
rect 8403 2040 8411 2074
rect 8445 2040 8453 2074
rect 8403 1915 8453 2040
rect 8489 2587 8497 2621
rect 8531 2587 8539 2621
rect 8489 2210 8539 2587
rect 8489 2176 8497 2210
rect 8531 2176 8539 2210
rect 8489 2142 8539 2176
rect 8489 2108 8497 2142
rect 8531 2108 8539 2142
rect 8489 2074 8539 2108
rect 8489 2040 8497 2074
rect 8531 2040 8539 2074
rect 8489 1915 8539 2040
rect 8575 2537 8625 2621
rect 8575 2503 8583 2537
rect 8617 2503 8625 2537
rect 8575 2210 8625 2503
rect 8575 2176 8583 2210
rect 8617 2176 8625 2210
rect 8575 2142 8625 2176
rect 8575 2108 8583 2142
rect 8617 2108 8625 2142
rect 8575 2074 8625 2108
rect 8575 2040 8583 2074
rect 8617 2040 8625 2074
rect 8575 1915 8625 2040
rect 8661 2587 8669 2621
rect 8703 2587 8711 2621
rect 8661 2210 8711 2587
rect 8661 2176 8669 2210
rect 8703 2176 8711 2210
rect 8661 2142 8711 2176
rect 8661 2108 8669 2142
rect 8703 2108 8711 2142
rect 8661 2074 8711 2108
rect 8661 2040 8669 2074
rect 8703 2040 8711 2074
rect 8661 1915 8711 2040
rect 8747 2537 8797 2621
rect 8747 2503 8755 2537
rect 8789 2503 8797 2537
rect 8747 2210 8797 2503
rect 8747 2176 8755 2210
rect 8789 2176 8797 2210
rect 8747 2142 8797 2176
rect 8747 2108 8755 2142
rect 8789 2108 8797 2142
rect 8747 2074 8797 2108
rect 8747 2040 8755 2074
rect 8789 2040 8797 2074
rect 8747 1915 8797 2040
rect 8833 2587 8841 2621
rect 8875 2587 8883 2621
rect 8833 2210 8883 2587
rect 8833 2176 8841 2210
rect 8875 2176 8883 2210
rect 8833 2142 8883 2176
rect 8833 2108 8841 2142
rect 8875 2108 8883 2142
rect 8833 2074 8883 2108
rect 8833 2040 8841 2074
rect 8875 2040 8883 2074
rect 8833 1915 8883 2040
rect 8919 2537 8969 2621
rect 8919 2503 8927 2537
rect 8961 2503 8969 2537
rect 8919 2210 8969 2503
rect 8919 2176 8927 2210
rect 8961 2176 8969 2210
rect 8919 2142 8969 2176
rect 8919 2108 8927 2142
rect 8961 2108 8969 2142
rect 8919 2074 8969 2108
rect 8919 2040 8927 2074
rect 8961 2040 8969 2074
rect 8919 1915 8969 2040
rect 9005 2587 9013 2621
rect 9047 2587 9055 2621
rect 9005 2210 9055 2587
rect 9005 2176 9013 2210
rect 9047 2176 9055 2210
rect 9005 2142 9055 2176
rect 9005 2108 9013 2142
rect 9047 2108 9055 2142
rect 9005 2074 9055 2108
rect 9005 2040 9013 2074
rect 9047 2040 9055 2074
rect 9005 1915 9055 2040
rect 9091 2537 9141 2621
rect 9091 2503 9099 2537
rect 9133 2503 9141 2537
rect 9091 2210 9141 2503
rect 9091 2176 9099 2210
rect 9133 2176 9141 2210
rect 9091 2142 9141 2176
rect 9091 2108 9099 2142
rect 9133 2108 9141 2142
rect 9091 2074 9141 2108
rect 9091 2040 9099 2074
rect 9133 2040 9141 2074
rect 9091 1915 9141 2040
rect 9177 2587 9185 2621
rect 9219 2587 9227 2621
rect 9177 2210 9227 2587
rect 9177 2176 9185 2210
rect 9219 2176 9227 2210
rect 9177 2142 9227 2176
rect 9177 2108 9185 2142
rect 9219 2108 9227 2142
rect 9177 2074 9227 2108
rect 9177 2040 9185 2074
rect 9219 2040 9227 2074
rect 9177 1915 9227 2040
rect 9263 2537 9313 2621
rect 9263 2503 9271 2537
rect 9305 2503 9313 2537
rect 9263 2210 9313 2503
rect 9263 2176 9271 2210
rect 9305 2176 9313 2210
rect 9263 2142 9313 2176
rect 9263 2108 9271 2142
rect 9305 2108 9313 2142
rect 9263 2074 9313 2108
rect 9263 2040 9271 2074
rect 9305 2040 9313 2074
rect 9263 1915 9313 2040
rect 9349 2587 9357 2621
rect 9391 2587 9399 2621
rect 9349 2210 9399 2587
rect 9349 2176 9357 2210
rect 9391 2176 9399 2210
rect 9349 2142 9399 2176
rect 9349 2108 9357 2142
rect 9391 2108 9399 2142
rect 9349 2074 9399 2108
rect 9349 2040 9357 2074
rect 9391 2040 9399 2074
rect 9349 1915 9399 2040
rect 9435 2537 9485 2621
rect 9435 2503 9443 2537
rect 9477 2503 9485 2537
rect 9435 2210 9485 2503
rect 9435 2176 9443 2210
rect 9477 2176 9485 2210
rect 9435 2142 9485 2176
rect 9435 2108 9443 2142
rect 9477 2108 9485 2142
rect 9435 2074 9485 2108
rect 9435 2040 9443 2074
rect 9477 2040 9485 2074
rect 9435 1915 9485 2040
rect 9521 2587 9529 2621
rect 9563 2587 9571 2621
rect 9521 2210 9571 2587
rect 9521 2176 9529 2210
rect 9563 2176 9571 2210
rect 9521 2142 9571 2176
rect 9521 2108 9529 2142
rect 9563 2108 9571 2142
rect 9521 2074 9571 2108
rect 9521 2040 9529 2074
rect 9563 2040 9571 2074
rect 9521 1915 9571 2040
rect 9607 2537 9657 2621
rect 9607 2503 9615 2537
rect 9649 2503 9657 2537
rect 9607 2210 9657 2503
rect 9607 2176 9615 2210
rect 9649 2176 9657 2210
rect 9607 2142 9657 2176
rect 9607 2108 9615 2142
rect 9649 2108 9657 2142
rect 9607 2074 9657 2108
rect 9607 2040 9615 2074
rect 9649 2040 9657 2074
rect 9607 1915 9657 2040
rect 9693 2587 9701 2621
rect 9735 2587 9743 2621
rect 9693 2210 9743 2587
rect 9693 2176 9701 2210
rect 9735 2176 9743 2210
rect 9693 2142 9743 2176
rect 9693 2108 9701 2142
rect 9735 2108 9743 2142
rect 9693 2074 9743 2108
rect 9693 2040 9701 2074
rect 9735 2040 9743 2074
rect 9693 1915 9743 2040
rect 9779 2537 9829 2621
rect 9779 2503 9787 2537
rect 9821 2503 9829 2537
rect 9779 2210 9829 2503
rect 9779 2176 9787 2210
rect 9821 2176 9829 2210
rect 9779 2142 9829 2176
rect 9779 2108 9787 2142
rect 9821 2108 9829 2142
rect 9779 2074 9829 2108
rect 9779 2040 9787 2074
rect 9821 2040 9829 2074
rect 9779 1915 9829 2040
rect 9865 2587 9873 2621
rect 9907 2587 9915 2621
rect 9865 2210 9915 2587
rect 9865 2176 9873 2210
rect 9907 2176 9915 2210
rect 9865 2142 9915 2176
rect 9865 2108 9873 2142
rect 9907 2108 9915 2142
rect 9865 2074 9915 2108
rect 9865 2040 9873 2074
rect 9907 2040 9915 2074
rect 9865 1915 9915 2040
rect 9951 2537 10001 2621
rect 9951 2503 9959 2537
rect 9993 2503 10001 2537
rect 9951 2210 10001 2503
rect 9951 2176 9959 2210
rect 9993 2176 10001 2210
rect 9951 2142 10001 2176
rect 9951 2108 9959 2142
rect 9993 2108 10001 2142
rect 9951 2074 10001 2108
rect 9951 2040 9959 2074
rect 9993 2040 10001 2074
rect 9951 1915 10001 2040
rect 10037 2587 10045 2621
rect 10079 2587 10087 2621
rect 10037 2210 10087 2587
rect 10037 2176 10045 2210
rect 10079 2176 10087 2210
rect 10037 2142 10087 2176
rect 10037 2108 10045 2142
rect 10079 2108 10087 2142
rect 10037 2074 10087 2108
rect 10037 2040 10045 2074
rect 10079 2040 10087 2074
rect 10037 1915 10087 2040
rect 10123 2537 10173 2621
rect 10123 2503 10131 2537
rect 10165 2503 10173 2537
rect 10123 2210 10173 2503
rect 10123 2176 10131 2210
rect 10165 2176 10173 2210
rect 10123 2142 10173 2176
rect 10123 2108 10131 2142
rect 10165 2108 10173 2142
rect 10123 2074 10173 2108
rect 10123 2040 10131 2074
rect 10165 2040 10173 2074
rect 10123 1915 10173 2040
rect 10209 2587 10217 2621
rect 10251 2587 10259 2621
rect 10209 2210 10259 2587
rect 10209 2176 10217 2210
rect 10251 2176 10259 2210
rect 10209 2142 10259 2176
rect 10209 2108 10217 2142
rect 10251 2108 10259 2142
rect 10209 2074 10259 2108
rect 10209 2040 10217 2074
rect 10251 2040 10259 2074
rect 10209 1915 10259 2040
rect 10295 2537 10345 2621
rect 10295 2503 10303 2537
rect 10337 2503 10345 2537
rect 10295 2210 10345 2503
rect 10295 2176 10303 2210
rect 10337 2176 10345 2210
rect 10295 2142 10345 2176
rect 10295 2108 10303 2142
rect 10337 2108 10345 2142
rect 10295 2074 10345 2108
rect 10295 2040 10303 2074
rect 10337 2040 10345 2074
rect 10295 1915 10345 2040
rect 10381 2587 10389 2621
rect 10423 2587 10431 2621
rect 10381 2210 10431 2587
rect 10381 2176 10389 2210
rect 10423 2176 10431 2210
rect 10381 2142 10431 2176
rect 10381 2108 10389 2142
rect 10423 2108 10431 2142
rect 10381 2074 10431 2108
rect 10381 2040 10389 2074
rect 10423 2040 10431 2074
rect 10381 1915 10431 2040
rect 10467 2537 10517 2621
rect 10467 2503 10475 2537
rect 10509 2503 10517 2537
rect 10467 2210 10517 2503
rect 10467 2176 10475 2210
rect 10509 2176 10517 2210
rect 10467 2142 10517 2176
rect 10467 2108 10475 2142
rect 10509 2108 10517 2142
rect 10467 2074 10517 2108
rect 10467 2040 10475 2074
rect 10509 2040 10517 2074
rect 10467 1915 10517 2040
rect 10553 2587 10561 2621
rect 10595 2587 10603 2621
rect 10553 2210 10603 2587
rect 10553 2176 10561 2210
rect 10595 2176 10603 2210
rect 10553 2142 10603 2176
rect 10553 2108 10561 2142
rect 10595 2108 10603 2142
rect 10553 2074 10603 2108
rect 10553 2040 10561 2074
rect 10595 2040 10603 2074
rect 10553 1915 10603 2040
rect 10639 2537 10689 2621
rect 10639 2503 10647 2537
rect 10681 2503 10689 2537
rect 10639 2210 10689 2503
rect 10639 2176 10647 2210
rect 10681 2176 10689 2210
rect 10639 2142 10689 2176
rect 10639 2108 10647 2142
rect 10681 2108 10689 2142
rect 10639 2074 10689 2108
rect 10639 2040 10647 2074
rect 10681 2040 10689 2074
rect 10639 1915 10689 2040
rect 10725 2587 10733 2621
rect 10767 2587 10775 2621
rect 10725 2210 10775 2587
rect 10725 2176 10733 2210
rect 10767 2176 10775 2210
rect 10725 2142 10775 2176
rect 10725 2108 10733 2142
rect 10767 2108 10775 2142
rect 10725 2074 10775 2108
rect 10725 2040 10733 2074
rect 10767 2040 10775 2074
rect 10725 1915 10775 2040
rect 10811 2537 10861 2621
rect 10811 2503 10819 2537
rect 10853 2503 10861 2537
rect 10811 2210 10861 2503
rect 10811 2176 10819 2210
rect 10853 2176 10861 2210
rect 10811 2142 10861 2176
rect 10811 2108 10819 2142
rect 10853 2108 10861 2142
rect 10811 2074 10861 2108
rect 10811 2040 10819 2074
rect 10853 2040 10861 2074
rect 10811 1915 10861 2040
rect 10897 2587 10905 2621
rect 10939 2587 10947 2621
rect 10897 2210 10947 2587
rect 10897 2176 10905 2210
rect 10939 2176 10947 2210
rect 10897 2142 10947 2176
rect 10897 2108 10905 2142
rect 10939 2108 10947 2142
rect 10897 2074 10947 2108
rect 10897 2040 10905 2074
rect 10939 2040 10947 2074
rect 10897 1915 10947 2040
rect 10983 2537 11033 2621
rect 10983 2503 10991 2537
rect 11025 2503 11033 2537
rect 10983 2210 11033 2503
rect 10983 2176 10991 2210
rect 11025 2176 11033 2210
rect 10983 2142 11033 2176
rect 10983 2108 10991 2142
rect 11025 2108 11033 2142
rect 10983 2074 11033 2108
rect 10983 2040 10991 2074
rect 11025 2040 11033 2074
rect 10983 1915 11033 2040
rect 11069 2587 11077 2621
rect 11111 2587 11119 2621
rect 11069 2210 11119 2587
rect 11069 2176 11077 2210
rect 11111 2176 11119 2210
rect 11069 2142 11119 2176
rect 11069 2108 11077 2142
rect 11111 2108 11119 2142
rect 11069 2074 11119 2108
rect 11069 2040 11077 2074
rect 11111 2040 11119 2074
rect 11069 1915 11119 2040
rect 11155 2537 11205 2621
rect 11155 2503 11163 2537
rect 11197 2503 11205 2537
rect 11155 2210 11205 2503
rect 11155 2176 11163 2210
rect 11197 2176 11205 2210
rect 11155 2142 11205 2176
rect 11155 2108 11163 2142
rect 11197 2108 11205 2142
rect 11155 2074 11205 2108
rect 11155 2040 11163 2074
rect 11197 2040 11205 2074
rect 11155 1915 11205 2040
rect 11241 2587 11249 2621
rect 11283 2587 11291 2621
rect 11241 2210 11291 2587
rect 11241 2176 11249 2210
rect 11283 2176 11291 2210
rect 11241 2142 11291 2176
rect 11241 2108 11249 2142
rect 11283 2108 11291 2142
rect 11241 2074 11291 2108
rect 11241 2040 11249 2074
rect 11283 2040 11291 2074
rect 11241 1915 11291 2040
rect 11327 2537 11377 2621
rect 11327 2503 11335 2537
rect 11369 2503 11377 2537
rect 11327 2210 11377 2503
rect 11327 2176 11335 2210
rect 11369 2176 11377 2210
rect 11327 2142 11377 2176
rect 11327 2108 11335 2142
rect 11369 2108 11377 2142
rect 11327 2074 11377 2108
rect 11327 2040 11335 2074
rect 11369 2040 11377 2074
rect 11327 1915 11377 2040
rect 5221 1865 5271 1915
rect 233 1781 283 1865
rect 233 1747 241 1781
rect 275 1747 283 1781
rect 233 1663 283 1747
rect 405 1781 455 1865
rect 405 1747 413 1781
rect 447 1747 455 1781
rect 405 1663 455 1747
rect 577 1781 627 1865
rect 577 1747 585 1781
rect 619 1747 627 1781
rect 577 1663 627 1747
rect 749 1781 799 1865
rect 749 1747 757 1781
rect 791 1747 799 1781
rect 749 1663 799 1747
rect 921 1781 971 1865
rect 921 1747 929 1781
rect 963 1747 971 1781
rect 921 1663 971 1747
rect 1093 1781 1143 1865
rect 1093 1747 1101 1781
rect 1135 1747 1143 1781
rect 1093 1663 1143 1747
rect 1265 1781 1315 1865
rect 1265 1747 1273 1781
rect 1307 1747 1315 1781
rect 1265 1663 1315 1747
rect 1437 1781 1487 1865
rect 1437 1747 1445 1781
rect 1479 1747 1487 1781
rect 1437 1663 1487 1747
rect 1609 1781 1659 1865
rect 1609 1747 1617 1781
rect 1651 1747 1659 1781
rect 1609 1663 1659 1747
rect 1781 1781 1831 1865
rect 1781 1747 1789 1781
rect 1823 1747 1831 1781
rect 1781 1663 1831 1747
rect 1953 1781 2003 1865
rect 1953 1747 1961 1781
rect 1995 1747 2003 1781
rect 1953 1663 2003 1747
rect 2125 1781 2175 1865
rect 2125 1747 2133 1781
rect 2167 1747 2175 1781
rect 2125 1663 2175 1747
rect 2641 1781 2691 1865
rect 2641 1747 2649 1781
rect 2683 1747 2691 1781
rect 2641 1663 2691 1747
rect 2813 1781 2863 1865
rect 2813 1747 2821 1781
rect 2855 1747 2863 1781
rect 2813 1663 2863 1747
rect 2985 1781 3035 1865
rect 2985 1747 2993 1781
rect 3027 1747 3035 1781
rect 2985 1663 3035 1747
rect 3157 1781 3207 1865
rect 3157 1747 3165 1781
rect 3199 1747 3207 1781
rect 3157 1663 3207 1747
rect 3329 1781 3379 1865
rect 3329 1747 3337 1781
rect 3371 1747 3379 1781
rect 3329 1663 3379 1747
rect 3501 1781 3551 1865
rect 3501 1747 3509 1781
rect 3543 1747 3551 1781
rect 3501 1663 3551 1747
rect 3931 1781 3981 1865
rect 3931 1747 3939 1781
rect 3973 1747 3981 1781
rect 3931 1454 3981 1747
rect 147 1361 197 1445
rect 147 1327 155 1361
rect 189 1327 197 1361
rect 147 1034 197 1327
rect 147 1000 155 1034
rect 189 1000 197 1034
rect 147 966 197 1000
rect 147 932 155 966
rect 189 932 197 966
rect 147 898 197 932
rect 147 864 155 898
rect 189 864 197 898
rect 147 739 197 864
rect 233 1411 241 1445
rect 275 1411 283 1445
rect 233 1034 283 1411
rect 233 1000 241 1034
rect 275 1000 283 1034
rect 233 966 283 1000
rect 233 932 241 966
rect 275 932 283 966
rect 233 898 283 932
rect 233 864 241 898
rect 275 864 283 898
rect 233 739 283 864
rect 319 1361 369 1445
rect 319 1327 327 1361
rect 361 1327 369 1361
rect 319 1034 369 1327
rect 319 1000 327 1034
rect 361 1000 369 1034
rect 319 966 369 1000
rect 319 932 327 966
rect 361 932 369 966
rect 319 898 369 932
rect 319 864 327 898
rect 361 864 369 898
rect 319 739 369 864
rect 405 1411 413 1445
rect 447 1411 455 1445
rect 405 1034 455 1411
rect 405 1000 413 1034
rect 447 1000 455 1034
rect 405 966 455 1000
rect 405 932 413 966
rect 447 932 455 966
rect 405 898 455 932
rect 405 864 413 898
rect 447 864 455 898
rect 405 739 455 864
rect 491 1361 541 1445
rect 491 1327 499 1361
rect 533 1327 541 1361
rect 491 1034 541 1327
rect 491 1000 499 1034
rect 533 1000 541 1034
rect 491 966 541 1000
rect 491 932 499 966
rect 533 932 541 966
rect 491 898 541 932
rect 491 864 499 898
rect 533 864 541 898
rect 491 739 541 864
rect 577 1411 585 1445
rect 619 1411 627 1445
rect 577 1034 627 1411
rect 577 1000 585 1034
rect 619 1000 627 1034
rect 577 966 627 1000
rect 577 932 585 966
rect 619 932 627 966
rect 577 898 627 932
rect 577 864 585 898
rect 619 864 627 898
rect 577 739 627 864
rect 663 1361 713 1445
rect 663 1327 671 1361
rect 705 1327 713 1361
rect 663 1034 713 1327
rect 663 1000 671 1034
rect 705 1000 713 1034
rect 663 966 713 1000
rect 663 932 671 966
rect 705 932 713 966
rect 663 898 713 932
rect 663 864 671 898
rect 705 864 713 898
rect 663 739 713 864
rect 749 1411 757 1445
rect 791 1411 799 1445
rect 749 1034 799 1411
rect 749 1000 757 1034
rect 791 1000 799 1034
rect 749 966 799 1000
rect 749 932 757 966
rect 791 932 799 966
rect 749 898 799 932
rect 749 864 757 898
rect 791 864 799 898
rect 749 739 799 864
rect 835 1361 885 1445
rect 835 1327 843 1361
rect 877 1327 885 1361
rect 835 1034 885 1327
rect 835 1000 843 1034
rect 877 1000 885 1034
rect 835 966 885 1000
rect 835 932 843 966
rect 877 932 885 966
rect 835 898 885 932
rect 835 864 843 898
rect 877 864 885 898
rect 835 739 885 864
rect 921 1411 929 1445
rect 963 1411 971 1445
rect 921 1034 971 1411
rect 921 1000 929 1034
rect 963 1000 971 1034
rect 921 966 971 1000
rect 921 932 929 966
rect 963 932 971 966
rect 921 898 971 932
rect 921 864 929 898
rect 963 864 971 898
rect 921 739 971 864
rect 1007 1361 1057 1445
rect 1007 1327 1015 1361
rect 1049 1327 1057 1361
rect 1007 1034 1057 1327
rect 1007 1000 1015 1034
rect 1049 1000 1057 1034
rect 1007 966 1057 1000
rect 1007 932 1015 966
rect 1049 932 1057 966
rect 1007 898 1057 932
rect 1007 864 1015 898
rect 1049 864 1057 898
rect 1007 739 1057 864
rect 1093 1411 1101 1445
rect 1135 1411 1143 1445
rect 1093 1034 1143 1411
rect 1093 1000 1101 1034
rect 1135 1000 1143 1034
rect 1093 966 1143 1000
rect 1093 932 1101 966
rect 1135 932 1143 966
rect 1093 898 1143 932
rect 1093 864 1101 898
rect 1135 864 1143 898
rect 1093 739 1143 864
rect 1179 1361 1229 1445
rect 1179 1327 1187 1361
rect 1221 1327 1229 1361
rect 1179 1034 1229 1327
rect 1179 1000 1187 1034
rect 1221 1000 1229 1034
rect 1179 966 1229 1000
rect 1179 932 1187 966
rect 1221 932 1229 966
rect 1179 898 1229 932
rect 1179 864 1187 898
rect 1221 864 1229 898
rect 1179 739 1229 864
rect 1265 1411 1273 1445
rect 1307 1411 1315 1445
rect 1265 1034 1315 1411
rect 1265 1000 1273 1034
rect 1307 1000 1315 1034
rect 1265 966 1315 1000
rect 1265 932 1273 966
rect 1307 932 1315 966
rect 1265 898 1315 932
rect 1265 864 1273 898
rect 1307 864 1315 898
rect 1265 739 1315 864
rect 1351 1361 1401 1445
rect 1351 1327 1359 1361
rect 1393 1327 1401 1361
rect 1351 1034 1401 1327
rect 1351 1000 1359 1034
rect 1393 1000 1401 1034
rect 1351 966 1401 1000
rect 1351 932 1359 966
rect 1393 932 1401 966
rect 1351 898 1401 932
rect 1351 864 1359 898
rect 1393 864 1401 898
rect 1351 739 1401 864
rect 1437 1411 1445 1445
rect 1479 1411 1487 1445
rect 1437 1034 1487 1411
rect 1437 1000 1445 1034
rect 1479 1000 1487 1034
rect 1437 966 1487 1000
rect 1437 932 1445 966
rect 1479 932 1487 966
rect 1437 898 1487 932
rect 1437 864 1445 898
rect 1479 864 1487 898
rect 1437 739 1487 864
rect 1523 1361 1573 1445
rect 1523 1327 1531 1361
rect 1565 1327 1573 1361
rect 1523 1034 1573 1327
rect 1523 1000 1531 1034
rect 1565 1000 1573 1034
rect 1523 966 1573 1000
rect 1523 932 1531 966
rect 1565 932 1573 966
rect 1523 898 1573 932
rect 1523 864 1531 898
rect 1565 864 1573 898
rect 1523 739 1573 864
rect 1609 1411 1617 1445
rect 1651 1411 1659 1445
rect 1609 1034 1659 1411
rect 1609 1000 1617 1034
rect 1651 1000 1659 1034
rect 1609 966 1659 1000
rect 1609 932 1617 966
rect 1651 932 1659 966
rect 1609 898 1659 932
rect 1609 864 1617 898
rect 1651 864 1659 898
rect 1609 739 1659 864
rect 1695 1361 1745 1445
rect 1695 1327 1703 1361
rect 1737 1327 1745 1361
rect 1695 1034 1745 1327
rect 1695 1000 1703 1034
rect 1737 1000 1745 1034
rect 1695 966 1745 1000
rect 1695 932 1703 966
rect 1737 932 1745 966
rect 1695 898 1745 932
rect 1695 864 1703 898
rect 1737 864 1745 898
rect 1695 739 1745 864
rect 1781 1411 1789 1445
rect 1823 1411 1831 1445
rect 1781 1034 1831 1411
rect 1781 1000 1789 1034
rect 1823 1000 1831 1034
rect 1781 966 1831 1000
rect 1781 932 1789 966
rect 1823 932 1831 966
rect 1781 898 1831 932
rect 1781 864 1789 898
rect 1823 864 1831 898
rect 1781 739 1831 864
rect 1867 1361 1917 1445
rect 1867 1327 1875 1361
rect 1909 1327 1917 1361
rect 1867 1034 1917 1327
rect 1867 1000 1875 1034
rect 1909 1000 1917 1034
rect 1867 966 1917 1000
rect 1867 932 1875 966
rect 1909 932 1917 966
rect 1867 898 1917 932
rect 1867 864 1875 898
rect 1909 864 1917 898
rect 1867 739 1917 864
rect 1953 1411 1961 1445
rect 1995 1411 2003 1445
rect 1953 1034 2003 1411
rect 1953 1000 1961 1034
rect 1995 1000 2003 1034
rect 1953 966 2003 1000
rect 1953 932 1961 966
rect 1995 932 2003 966
rect 1953 898 2003 932
rect 1953 864 1961 898
rect 1995 864 2003 898
rect 1953 739 2003 864
rect 2039 1361 2089 1445
rect 2039 1327 2047 1361
rect 2081 1327 2089 1361
rect 2039 1034 2089 1327
rect 2039 1000 2047 1034
rect 2081 1000 2089 1034
rect 2039 966 2089 1000
rect 2039 932 2047 966
rect 2081 932 2089 966
rect 2039 898 2089 932
rect 2039 864 2047 898
rect 2081 864 2089 898
rect 2039 739 2089 864
rect 2125 1411 2133 1445
rect 2167 1411 2175 1445
rect 2125 1034 2175 1411
rect 2125 1000 2133 1034
rect 2167 1000 2175 1034
rect 2125 966 2175 1000
rect 2125 932 2133 966
rect 2167 932 2175 966
rect 2125 898 2175 932
rect 2125 864 2133 898
rect 2167 864 2175 898
rect 2125 739 2175 864
rect 2211 1361 2261 1445
rect 2211 1327 2219 1361
rect 2253 1327 2261 1361
rect 2211 1034 2261 1327
rect 2211 1000 2219 1034
rect 2253 1000 2261 1034
rect 2211 966 2261 1000
rect 2211 932 2219 966
rect 2253 932 2261 966
rect 2211 898 2261 932
rect 2211 864 2219 898
rect 2253 864 2261 898
rect 2211 739 2261 864
rect 2555 1361 2605 1445
rect 2555 1327 2563 1361
rect 2597 1327 2605 1361
rect 2555 1034 2605 1327
rect 2555 1000 2563 1034
rect 2597 1000 2605 1034
rect 2555 966 2605 1000
rect 2555 932 2563 966
rect 2597 932 2605 966
rect 2555 898 2605 932
rect 2555 864 2563 898
rect 2597 864 2605 898
rect 2555 739 2605 864
rect 2641 1411 2649 1445
rect 2683 1411 2691 1445
rect 2641 1034 2691 1411
rect 2641 1000 2649 1034
rect 2683 1000 2691 1034
rect 2641 966 2691 1000
rect 2641 932 2649 966
rect 2683 932 2691 966
rect 2641 898 2691 932
rect 2641 864 2649 898
rect 2683 864 2691 898
rect 2641 739 2691 864
rect 2727 1361 2777 1445
rect 2727 1327 2735 1361
rect 2769 1327 2777 1361
rect 2727 1034 2777 1327
rect 2727 1000 2735 1034
rect 2769 1000 2777 1034
rect 2727 966 2777 1000
rect 2727 932 2735 966
rect 2769 932 2777 966
rect 2727 898 2777 932
rect 2727 864 2735 898
rect 2769 864 2777 898
rect 2727 739 2777 864
rect 2813 1411 2821 1445
rect 2855 1411 2863 1445
rect 2813 1034 2863 1411
rect 2813 1000 2821 1034
rect 2855 1000 2863 1034
rect 2813 966 2863 1000
rect 2813 932 2821 966
rect 2855 932 2863 966
rect 2813 898 2863 932
rect 2813 864 2821 898
rect 2855 864 2863 898
rect 2813 739 2863 864
rect 2899 1361 2949 1445
rect 2899 1327 2907 1361
rect 2941 1327 2949 1361
rect 2899 1034 2949 1327
rect 2899 1000 2907 1034
rect 2941 1000 2949 1034
rect 2899 966 2949 1000
rect 2899 932 2907 966
rect 2941 932 2949 966
rect 2899 898 2949 932
rect 2899 864 2907 898
rect 2941 864 2949 898
rect 2899 739 2949 864
rect 2985 1411 2993 1445
rect 3027 1411 3035 1445
rect 2985 1034 3035 1411
rect 2985 1000 2993 1034
rect 3027 1000 3035 1034
rect 2985 966 3035 1000
rect 2985 932 2993 966
rect 3027 932 3035 966
rect 2985 898 3035 932
rect 2985 864 2993 898
rect 3027 864 3035 898
rect 2985 739 3035 864
rect 3071 1361 3121 1445
rect 3071 1327 3079 1361
rect 3113 1327 3121 1361
rect 3071 1034 3121 1327
rect 3071 1000 3079 1034
rect 3113 1000 3121 1034
rect 3071 966 3121 1000
rect 3071 932 3079 966
rect 3113 932 3121 966
rect 3071 898 3121 932
rect 3071 864 3079 898
rect 3113 864 3121 898
rect 3071 739 3121 864
rect 3157 1411 3165 1445
rect 3199 1411 3207 1445
rect 3157 1034 3207 1411
rect 3157 1000 3165 1034
rect 3199 1000 3207 1034
rect 3157 966 3207 1000
rect 3157 932 3165 966
rect 3199 932 3207 966
rect 3157 898 3207 932
rect 3157 864 3165 898
rect 3199 864 3207 898
rect 3157 739 3207 864
rect 3243 1361 3293 1445
rect 3243 1327 3251 1361
rect 3285 1327 3293 1361
rect 3243 1034 3293 1327
rect 3243 1000 3251 1034
rect 3285 1000 3293 1034
rect 3243 966 3293 1000
rect 3243 932 3251 966
rect 3285 932 3293 966
rect 3243 898 3293 932
rect 3243 864 3251 898
rect 3285 864 3293 898
rect 3243 739 3293 864
rect 3329 1411 3337 1445
rect 3371 1411 3379 1445
rect 3329 1034 3379 1411
rect 3329 1000 3337 1034
rect 3371 1000 3379 1034
rect 3329 966 3379 1000
rect 3329 932 3337 966
rect 3371 932 3379 966
rect 3329 898 3379 932
rect 3329 864 3337 898
rect 3371 864 3379 898
rect 3329 739 3379 864
rect 3415 1361 3465 1445
rect 3415 1327 3423 1361
rect 3457 1327 3465 1361
rect 3415 1034 3465 1327
rect 3415 1000 3423 1034
rect 3457 1000 3465 1034
rect 3415 966 3465 1000
rect 3415 932 3423 966
rect 3457 932 3465 966
rect 3415 898 3465 932
rect 3415 864 3423 898
rect 3457 864 3465 898
rect 3415 739 3465 864
rect 3501 1411 3509 1445
rect 3543 1411 3551 1445
rect 3501 1034 3551 1411
rect 3501 1000 3509 1034
rect 3543 1000 3551 1034
rect 3501 966 3551 1000
rect 3501 932 3509 966
rect 3543 932 3551 966
rect 3501 898 3551 932
rect 3501 864 3509 898
rect 3543 864 3551 898
rect 3501 739 3551 864
rect 3587 1361 3637 1445
rect 3587 1327 3595 1361
rect 3629 1327 3637 1361
rect 3587 1034 3637 1327
rect 3931 1420 3939 1454
rect 3973 1420 3981 1454
rect 3931 1386 3981 1420
rect 3931 1352 3939 1386
rect 3973 1352 3981 1386
rect 3931 1318 3981 1352
rect 3931 1284 3939 1318
rect 3973 1284 3981 1318
rect 3931 1159 3981 1284
rect 4017 1831 4025 1865
rect 4059 1831 4067 1865
rect 4017 1454 4067 1831
rect 4017 1420 4025 1454
rect 4059 1420 4067 1454
rect 4017 1386 4067 1420
rect 4017 1352 4025 1386
rect 4059 1352 4067 1386
rect 4017 1318 4067 1352
rect 4017 1284 4025 1318
rect 4059 1284 4067 1318
rect 4017 1159 4067 1284
rect 4103 1781 4153 1865
rect 4103 1747 4111 1781
rect 4145 1747 4153 1781
rect 4103 1454 4153 1747
rect 4103 1420 4111 1454
rect 4145 1420 4153 1454
rect 4103 1386 4153 1420
rect 4103 1352 4111 1386
rect 4145 1352 4153 1386
rect 4103 1318 4153 1352
rect 4103 1284 4111 1318
rect 4145 1284 4153 1318
rect 4103 1159 4153 1284
rect 4189 1831 4197 1865
rect 4231 1831 4239 1865
rect 4189 1454 4239 1831
rect 4189 1420 4197 1454
rect 4231 1420 4239 1454
rect 4189 1386 4239 1420
rect 4189 1352 4197 1386
rect 4231 1352 4239 1386
rect 4189 1318 4239 1352
rect 4189 1284 4197 1318
rect 4231 1284 4239 1318
rect 4189 1159 4239 1284
rect 4275 1781 4325 1865
rect 4275 1747 4283 1781
rect 4317 1747 4325 1781
rect 4275 1454 4325 1747
rect 4275 1420 4283 1454
rect 4317 1420 4325 1454
rect 4275 1386 4325 1420
rect 4275 1352 4283 1386
rect 4317 1352 4325 1386
rect 4275 1318 4325 1352
rect 4275 1284 4283 1318
rect 4317 1284 4325 1318
rect 4275 1159 4325 1284
rect 4361 1831 4369 1865
rect 4403 1831 4411 1865
rect 4361 1454 4411 1831
rect 4361 1420 4369 1454
rect 4403 1420 4411 1454
rect 4361 1386 4411 1420
rect 4361 1352 4369 1386
rect 4403 1352 4411 1386
rect 4361 1318 4411 1352
rect 4361 1284 4369 1318
rect 4403 1284 4411 1318
rect 4361 1159 4411 1284
rect 4447 1781 4497 1865
rect 4447 1747 4455 1781
rect 4489 1747 4497 1781
rect 4447 1454 4497 1747
rect 4447 1420 4455 1454
rect 4489 1420 4497 1454
rect 4447 1386 4497 1420
rect 4447 1352 4455 1386
rect 4489 1352 4497 1386
rect 4447 1318 4497 1352
rect 4447 1284 4455 1318
rect 4489 1284 4497 1318
rect 4447 1159 4497 1284
rect 4533 1831 4541 1865
rect 4575 1831 4583 1865
rect 4533 1454 4583 1831
rect 4533 1420 4541 1454
rect 4575 1420 4583 1454
rect 4533 1386 4583 1420
rect 4533 1352 4541 1386
rect 4575 1352 4583 1386
rect 4533 1318 4583 1352
rect 4533 1284 4541 1318
rect 4575 1284 4583 1318
rect 4533 1159 4583 1284
rect 4619 1781 4669 1865
rect 4619 1747 4627 1781
rect 4661 1747 4669 1781
rect 4619 1454 4669 1747
rect 4619 1420 4627 1454
rect 4661 1420 4669 1454
rect 4619 1386 4669 1420
rect 4619 1352 4627 1386
rect 4661 1352 4669 1386
rect 4619 1318 4669 1352
rect 4619 1284 4627 1318
rect 4661 1284 4669 1318
rect 4619 1159 4669 1284
rect 4705 1831 4713 1865
rect 4747 1831 4755 1865
rect 4705 1454 4755 1831
rect 4705 1420 4713 1454
rect 4747 1420 4755 1454
rect 4705 1386 4755 1420
rect 4705 1352 4713 1386
rect 4747 1352 4755 1386
rect 4705 1318 4755 1352
rect 4705 1284 4713 1318
rect 4747 1284 4755 1318
rect 4705 1159 4755 1284
rect 4791 1781 4841 1865
rect 4791 1747 4799 1781
rect 4833 1747 4841 1781
rect 4791 1454 4841 1747
rect 4791 1420 4799 1454
rect 4833 1420 4841 1454
rect 4791 1386 4841 1420
rect 4791 1352 4799 1386
rect 4833 1352 4841 1386
rect 4791 1318 4841 1352
rect 4791 1284 4799 1318
rect 4833 1284 4841 1318
rect 4791 1159 4841 1284
rect 4877 1831 4885 1865
rect 4919 1831 4927 1865
rect 4877 1454 4927 1831
rect 4877 1420 4885 1454
rect 4919 1420 4927 1454
rect 4877 1386 4927 1420
rect 4877 1352 4885 1386
rect 4919 1352 4927 1386
rect 4877 1318 4927 1352
rect 4877 1284 4885 1318
rect 4919 1284 4927 1318
rect 4877 1159 4927 1284
rect 4963 1781 5013 1865
rect 5221 1831 5229 1865
rect 5263 1831 5271 1865
rect 4963 1747 4971 1781
rect 5005 1747 5013 1781
rect 4963 1454 5013 1747
rect 4963 1420 4971 1454
rect 5005 1420 5013 1454
rect 4963 1386 5013 1420
rect 4963 1352 4971 1386
rect 5005 1352 5013 1386
rect 4963 1318 5013 1352
rect 4963 1284 4971 1318
rect 5005 1284 5013 1318
rect 4963 1159 5013 1284
rect 5307 1781 5357 1865
rect 5307 1747 5315 1781
rect 5349 1747 5357 1781
rect 5307 1454 5357 1747
rect 5307 1420 5315 1454
rect 5349 1420 5357 1454
rect 5307 1386 5357 1420
rect 5307 1352 5315 1386
rect 5349 1352 5357 1386
rect 5307 1318 5357 1352
rect 5307 1284 5315 1318
rect 5349 1284 5357 1318
rect 5307 1159 5357 1284
rect 5393 1831 5401 1865
rect 5435 1831 5443 1865
rect 5393 1454 5443 1831
rect 5393 1420 5401 1454
rect 5435 1420 5443 1454
rect 5393 1386 5443 1420
rect 5393 1352 5401 1386
rect 5435 1352 5443 1386
rect 5393 1318 5443 1352
rect 5393 1284 5401 1318
rect 5435 1284 5443 1318
rect 5393 1159 5443 1284
rect 5479 1781 5529 1865
rect 5479 1747 5487 1781
rect 5521 1747 5529 1781
rect 5479 1454 5529 1747
rect 5479 1420 5487 1454
rect 5521 1420 5529 1454
rect 5479 1386 5529 1420
rect 5479 1352 5487 1386
rect 5521 1352 5529 1386
rect 5479 1318 5529 1352
rect 5479 1284 5487 1318
rect 5521 1284 5529 1318
rect 5479 1159 5529 1284
rect 5565 1831 5573 1865
rect 5607 1831 5615 1865
rect 5565 1454 5615 1831
rect 5565 1420 5573 1454
rect 5607 1420 5615 1454
rect 5565 1386 5615 1420
rect 5565 1352 5573 1386
rect 5607 1352 5615 1386
rect 5565 1318 5615 1352
rect 5565 1284 5573 1318
rect 5607 1284 5615 1318
rect 5565 1159 5615 1284
rect 5651 1781 5701 1865
rect 5651 1747 5659 1781
rect 5693 1747 5701 1781
rect 5651 1454 5701 1747
rect 5651 1420 5659 1454
rect 5693 1420 5701 1454
rect 5651 1386 5701 1420
rect 5651 1352 5659 1386
rect 5693 1352 5701 1386
rect 5651 1318 5701 1352
rect 5651 1284 5659 1318
rect 5693 1284 5701 1318
rect 5651 1159 5701 1284
rect 5737 1831 5745 1865
rect 5779 1831 5787 1865
rect 5737 1454 5787 1831
rect 5737 1420 5745 1454
rect 5779 1420 5787 1454
rect 5737 1386 5787 1420
rect 5737 1352 5745 1386
rect 5779 1352 5787 1386
rect 5737 1318 5787 1352
rect 5737 1284 5745 1318
rect 5779 1284 5787 1318
rect 5737 1159 5787 1284
rect 5823 1781 5873 1865
rect 5823 1747 5831 1781
rect 5865 1747 5873 1781
rect 5823 1454 5873 1747
rect 6253 1781 6303 1865
rect 6253 1747 6261 1781
rect 6295 1747 6303 1781
rect 6253 1663 6303 1747
rect 6769 1781 6819 1865
rect 6769 1747 6777 1781
rect 6811 1747 6819 1781
rect 6769 1663 6819 1747
rect 7285 1781 7335 1865
rect 7285 1747 7293 1781
rect 7327 1747 7335 1781
rect 7285 1663 7335 1747
rect 7457 1781 7507 1865
rect 7457 1747 7465 1781
rect 7499 1747 7507 1781
rect 7457 1663 7507 1747
rect 7629 1781 7679 1865
rect 7629 1747 7637 1781
rect 7671 1747 7679 1781
rect 7629 1663 7679 1747
rect 7801 1781 7851 1865
rect 7801 1747 7809 1781
rect 7843 1747 7851 1781
rect 7801 1663 7851 1747
rect 7973 1781 8023 1865
rect 7973 1747 7981 1781
rect 8015 1747 8023 1781
rect 7973 1663 8023 1747
rect 8145 1781 8195 1865
rect 8145 1747 8153 1781
rect 8187 1747 8195 1781
rect 8145 1663 8195 1747
rect 8317 1781 8367 1865
rect 8317 1747 8325 1781
rect 8359 1747 8367 1781
rect 8317 1663 8367 1747
rect 8489 1781 8539 1865
rect 8489 1747 8497 1781
rect 8531 1747 8539 1781
rect 8489 1663 8539 1747
rect 8661 1781 8711 1865
rect 8661 1747 8669 1781
rect 8703 1747 8711 1781
rect 8661 1663 8711 1747
rect 8833 1781 8883 1865
rect 8833 1747 8841 1781
rect 8875 1747 8883 1781
rect 8833 1663 8883 1747
rect 9005 1781 9055 1865
rect 9005 1747 9013 1781
rect 9047 1747 9055 1781
rect 9005 1663 9055 1747
rect 9177 1781 9227 1865
rect 9177 1747 9185 1781
rect 9219 1747 9227 1781
rect 9177 1663 9227 1747
rect 9349 1781 9399 1865
rect 9349 1747 9357 1781
rect 9391 1747 9399 1781
rect 9349 1663 9399 1747
rect 9521 1781 9571 1865
rect 9521 1747 9529 1781
rect 9563 1747 9571 1781
rect 9521 1663 9571 1747
rect 9693 1781 9743 1865
rect 9693 1747 9701 1781
rect 9735 1747 9743 1781
rect 9693 1663 9743 1747
rect 9865 1781 9915 1865
rect 9865 1747 9873 1781
rect 9907 1747 9915 1781
rect 9865 1663 9915 1747
rect 10037 1781 10087 1865
rect 10037 1747 10045 1781
rect 10079 1747 10087 1781
rect 10037 1663 10087 1747
rect 10209 1781 10259 1865
rect 10209 1747 10217 1781
rect 10251 1747 10259 1781
rect 10209 1663 10259 1747
rect 10381 1781 10431 1865
rect 10381 1747 10389 1781
rect 10423 1747 10431 1781
rect 10381 1663 10431 1747
rect 10553 1781 10603 1865
rect 10553 1747 10561 1781
rect 10595 1747 10603 1781
rect 10553 1663 10603 1747
rect 10725 1781 10775 1865
rect 10725 1747 10733 1781
rect 10767 1747 10775 1781
rect 10725 1663 10775 1747
rect 10897 1781 10947 1865
rect 10897 1747 10905 1781
rect 10939 1747 10947 1781
rect 10897 1663 10947 1747
rect 11069 1781 11119 1865
rect 11069 1747 11077 1781
rect 11111 1747 11119 1781
rect 11069 1663 11119 1747
rect 11241 1781 11291 1865
rect 11241 1747 11249 1781
rect 11283 1747 11291 1781
rect 11241 1663 11291 1747
rect 5823 1420 5831 1454
rect 5865 1420 5873 1454
rect 5823 1386 5873 1420
rect 5823 1352 5831 1386
rect 5865 1352 5873 1386
rect 5823 1318 5873 1352
rect 5823 1284 5831 1318
rect 5865 1284 5873 1318
rect 5823 1159 5873 1284
rect 6167 1488 6217 1613
rect 6167 1454 6175 1488
rect 6209 1454 6217 1488
rect 6167 1420 6217 1454
rect 6167 1386 6175 1420
rect 6209 1386 6217 1420
rect 6167 1352 6217 1386
rect 6167 1318 6175 1352
rect 6209 1318 6217 1352
rect 3587 1000 3595 1034
rect 3629 1000 3637 1034
rect 3587 966 3637 1000
rect 3587 932 3595 966
rect 3629 932 3637 966
rect 3587 898 3637 932
rect 4017 1025 4067 1109
rect 4017 991 4025 1025
rect 4059 991 4067 1025
rect 4017 907 4067 991
rect 4189 1025 4239 1109
rect 4189 991 4197 1025
rect 4231 991 4239 1025
rect 4189 907 4239 991
rect 4361 1025 4411 1109
rect 4361 991 4369 1025
rect 4403 991 4411 1025
rect 4361 907 4411 991
rect 4533 1025 4583 1109
rect 4533 991 4541 1025
rect 4575 991 4583 1025
rect 4533 907 4583 991
rect 4705 1025 4755 1109
rect 4705 991 4713 1025
rect 4747 991 4755 1025
rect 4705 907 4755 991
rect 4877 1025 4927 1109
rect 4877 991 4885 1025
rect 4919 991 4927 1025
rect 4877 907 4927 991
rect 5393 1025 5443 1109
rect 5393 991 5401 1025
rect 5435 991 5443 1025
rect 5393 907 5443 991
rect 5565 1025 5615 1109
rect 5565 991 5573 1025
rect 5607 991 5615 1025
rect 5565 907 5615 991
rect 5737 1025 5787 1109
rect 5737 991 5745 1025
rect 5779 991 5787 1025
rect 5737 907 5787 991
rect 6167 1025 6217 1318
rect 6167 991 6175 1025
rect 6209 991 6217 1025
rect 6167 907 6217 991
rect 6253 1488 6303 1613
rect 6253 1454 6261 1488
rect 6295 1454 6303 1488
rect 6253 1420 6303 1454
rect 6253 1386 6261 1420
rect 6295 1386 6303 1420
rect 6253 1352 6303 1386
rect 6253 1318 6261 1352
rect 6295 1318 6303 1352
rect 6253 941 6303 1318
rect 6253 907 6261 941
rect 6295 907 6303 941
rect 6339 1488 6389 1613
rect 6339 1454 6347 1488
rect 6381 1454 6389 1488
rect 6339 1420 6389 1454
rect 6339 1386 6347 1420
rect 6381 1386 6389 1420
rect 6339 1352 6389 1386
rect 6339 1318 6347 1352
rect 6381 1318 6389 1352
rect 6339 1025 6389 1318
rect 6769 1361 6819 1445
rect 6769 1327 6777 1361
rect 6811 1327 6819 1361
rect 6769 1243 6819 1327
rect 7199 1361 7249 1445
rect 7199 1327 7207 1361
rect 7241 1327 7249 1361
rect 6339 991 6347 1025
rect 6381 991 6389 1025
rect 6339 907 6389 991
rect 7199 1034 7249 1327
rect 7199 1000 7207 1034
rect 7241 1000 7249 1034
rect 7199 966 7249 1000
rect 7199 932 7207 966
rect 7241 932 7249 966
rect 3587 864 3595 898
rect 3629 864 3637 898
rect 3587 739 3637 864
rect 7199 898 7249 932
rect 7199 864 7207 898
rect 7241 864 7249 898
rect 7199 739 7249 864
rect 7285 1411 7293 1445
rect 7327 1411 7335 1445
rect 7285 1034 7335 1411
rect 7285 1000 7293 1034
rect 7327 1000 7335 1034
rect 7285 966 7335 1000
rect 7285 932 7293 966
rect 7327 932 7335 966
rect 7285 898 7335 932
rect 7285 864 7293 898
rect 7327 864 7335 898
rect 7285 739 7335 864
rect 7371 1361 7421 1445
rect 7371 1327 7379 1361
rect 7413 1327 7421 1361
rect 7371 1034 7421 1327
rect 7371 1000 7379 1034
rect 7413 1000 7421 1034
rect 7371 966 7421 1000
rect 7371 932 7379 966
rect 7413 932 7421 966
rect 7371 898 7421 932
rect 7371 864 7379 898
rect 7413 864 7421 898
rect 7371 739 7421 864
rect 7457 1411 7465 1445
rect 7499 1411 7507 1445
rect 7457 1034 7507 1411
rect 7457 1000 7465 1034
rect 7499 1000 7507 1034
rect 7457 966 7507 1000
rect 7457 932 7465 966
rect 7499 932 7507 966
rect 7457 898 7507 932
rect 7457 864 7465 898
rect 7499 864 7507 898
rect 7457 739 7507 864
rect 7543 1361 7593 1445
rect 7543 1327 7551 1361
rect 7585 1327 7593 1361
rect 7543 1034 7593 1327
rect 7543 1000 7551 1034
rect 7585 1000 7593 1034
rect 7543 966 7593 1000
rect 7543 932 7551 966
rect 7585 932 7593 966
rect 7543 898 7593 932
rect 7543 864 7551 898
rect 7585 864 7593 898
rect 7543 739 7593 864
rect 7629 1411 7637 1445
rect 7671 1411 7679 1445
rect 7629 1034 7679 1411
rect 7629 1000 7637 1034
rect 7671 1000 7679 1034
rect 7629 966 7679 1000
rect 7629 932 7637 966
rect 7671 932 7679 966
rect 7629 898 7679 932
rect 7629 864 7637 898
rect 7671 864 7679 898
rect 7629 739 7679 864
rect 7715 1361 7765 1445
rect 7715 1327 7723 1361
rect 7757 1327 7765 1361
rect 7715 1034 7765 1327
rect 7715 1000 7723 1034
rect 7757 1000 7765 1034
rect 7715 966 7765 1000
rect 7715 932 7723 966
rect 7757 932 7765 966
rect 7715 898 7765 932
rect 7715 864 7723 898
rect 7757 864 7765 898
rect 7715 739 7765 864
rect 7801 1411 7809 1445
rect 7843 1411 7851 1445
rect 7801 1034 7851 1411
rect 7801 1000 7809 1034
rect 7843 1000 7851 1034
rect 7801 966 7851 1000
rect 7801 932 7809 966
rect 7843 932 7851 966
rect 7801 898 7851 932
rect 7801 864 7809 898
rect 7843 864 7851 898
rect 7801 739 7851 864
rect 7887 1361 7937 1445
rect 7887 1327 7895 1361
rect 7929 1327 7937 1361
rect 7887 1034 7937 1327
rect 7887 1000 7895 1034
rect 7929 1000 7937 1034
rect 7887 966 7937 1000
rect 7887 932 7895 966
rect 7929 932 7937 966
rect 7887 898 7937 932
rect 7887 864 7895 898
rect 7929 864 7937 898
rect 7887 739 7937 864
rect 7973 1411 7981 1445
rect 8015 1411 8023 1445
rect 7973 1034 8023 1411
rect 7973 1000 7981 1034
rect 8015 1000 8023 1034
rect 7973 966 8023 1000
rect 7973 932 7981 966
rect 8015 932 8023 966
rect 7973 898 8023 932
rect 7973 864 7981 898
rect 8015 864 8023 898
rect 7973 739 8023 864
rect 8059 1361 8109 1445
rect 8059 1327 8067 1361
rect 8101 1327 8109 1361
rect 8059 1034 8109 1327
rect 8059 1000 8067 1034
rect 8101 1000 8109 1034
rect 8059 966 8109 1000
rect 8059 932 8067 966
rect 8101 932 8109 966
rect 8059 898 8109 932
rect 8059 864 8067 898
rect 8101 864 8109 898
rect 8059 739 8109 864
rect 8145 1411 8153 1445
rect 8187 1411 8195 1445
rect 8145 1034 8195 1411
rect 8145 1000 8153 1034
rect 8187 1000 8195 1034
rect 8145 966 8195 1000
rect 8145 932 8153 966
rect 8187 932 8195 966
rect 8145 898 8195 932
rect 8145 864 8153 898
rect 8187 864 8195 898
rect 8145 739 8195 864
rect 8231 1361 8281 1445
rect 8231 1327 8239 1361
rect 8273 1327 8281 1361
rect 8231 1034 8281 1327
rect 8231 1000 8239 1034
rect 8273 1000 8281 1034
rect 8231 966 8281 1000
rect 8231 932 8239 966
rect 8273 932 8281 966
rect 8231 898 8281 932
rect 8231 864 8239 898
rect 8273 864 8281 898
rect 8231 739 8281 864
rect 8317 1411 8325 1445
rect 8359 1411 8367 1445
rect 8317 1034 8367 1411
rect 8317 1000 8325 1034
rect 8359 1000 8367 1034
rect 8317 966 8367 1000
rect 8317 932 8325 966
rect 8359 932 8367 966
rect 8317 898 8367 932
rect 8317 864 8325 898
rect 8359 864 8367 898
rect 8317 739 8367 864
rect 8403 1361 8453 1445
rect 8403 1327 8411 1361
rect 8445 1327 8453 1361
rect 8403 1034 8453 1327
rect 8403 1000 8411 1034
rect 8445 1000 8453 1034
rect 8403 966 8453 1000
rect 8403 932 8411 966
rect 8445 932 8453 966
rect 8403 898 8453 932
rect 8403 864 8411 898
rect 8445 864 8453 898
rect 8403 739 8453 864
rect 8489 1411 8497 1445
rect 8531 1411 8539 1445
rect 8489 1034 8539 1411
rect 8489 1000 8497 1034
rect 8531 1000 8539 1034
rect 8489 966 8539 1000
rect 8489 932 8497 966
rect 8531 932 8539 966
rect 8489 898 8539 932
rect 8489 864 8497 898
rect 8531 864 8539 898
rect 8489 739 8539 864
rect 8575 1361 8625 1445
rect 8575 1327 8583 1361
rect 8617 1327 8625 1361
rect 8575 1034 8625 1327
rect 8575 1000 8583 1034
rect 8617 1000 8625 1034
rect 8575 966 8625 1000
rect 8575 932 8583 966
rect 8617 932 8625 966
rect 8575 898 8625 932
rect 8575 864 8583 898
rect 8617 864 8625 898
rect 8575 739 8625 864
rect 8661 1411 8669 1445
rect 8703 1411 8711 1445
rect 8661 1034 8711 1411
rect 8661 1000 8669 1034
rect 8703 1000 8711 1034
rect 8661 966 8711 1000
rect 8661 932 8669 966
rect 8703 932 8711 966
rect 8661 898 8711 932
rect 8661 864 8669 898
rect 8703 864 8711 898
rect 8661 739 8711 864
rect 8747 1361 8797 1445
rect 8747 1327 8755 1361
rect 8789 1327 8797 1361
rect 8747 1034 8797 1327
rect 8747 1000 8755 1034
rect 8789 1000 8797 1034
rect 8747 966 8797 1000
rect 8747 932 8755 966
rect 8789 932 8797 966
rect 8747 898 8797 932
rect 8747 864 8755 898
rect 8789 864 8797 898
rect 8747 739 8797 864
rect 8833 1411 8841 1445
rect 8875 1411 8883 1445
rect 8833 1034 8883 1411
rect 8833 1000 8841 1034
rect 8875 1000 8883 1034
rect 8833 966 8883 1000
rect 8833 932 8841 966
rect 8875 932 8883 966
rect 8833 898 8883 932
rect 8833 864 8841 898
rect 8875 864 8883 898
rect 8833 739 8883 864
rect 8919 1361 8969 1445
rect 8919 1327 8927 1361
rect 8961 1327 8969 1361
rect 8919 1034 8969 1327
rect 8919 1000 8927 1034
rect 8961 1000 8969 1034
rect 8919 966 8969 1000
rect 8919 932 8927 966
rect 8961 932 8969 966
rect 8919 898 8969 932
rect 8919 864 8927 898
rect 8961 864 8969 898
rect 8919 739 8969 864
rect 9005 1411 9013 1445
rect 9047 1411 9055 1445
rect 9005 1034 9055 1411
rect 9005 1000 9013 1034
rect 9047 1000 9055 1034
rect 9005 966 9055 1000
rect 9005 932 9013 966
rect 9047 932 9055 966
rect 9005 898 9055 932
rect 9005 864 9013 898
rect 9047 864 9055 898
rect 9005 739 9055 864
rect 9091 1361 9141 1445
rect 9091 1327 9099 1361
rect 9133 1327 9141 1361
rect 9091 1034 9141 1327
rect 9091 1000 9099 1034
rect 9133 1000 9141 1034
rect 9091 966 9141 1000
rect 9091 932 9099 966
rect 9133 932 9141 966
rect 9091 898 9141 932
rect 9091 864 9099 898
rect 9133 864 9141 898
rect 9091 739 9141 864
rect 9177 1411 9185 1445
rect 9219 1411 9227 1445
rect 9177 1034 9227 1411
rect 9177 1000 9185 1034
rect 9219 1000 9227 1034
rect 9177 966 9227 1000
rect 9177 932 9185 966
rect 9219 932 9227 966
rect 9177 898 9227 932
rect 9177 864 9185 898
rect 9219 864 9227 898
rect 9177 739 9227 864
rect 9263 1361 9313 1445
rect 9263 1327 9271 1361
rect 9305 1327 9313 1361
rect 9263 1034 9313 1327
rect 9263 1000 9271 1034
rect 9305 1000 9313 1034
rect 9263 966 9313 1000
rect 9263 932 9271 966
rect 9305 932 9313 966
rect 9263 898 9313 932
rect 9263 864 9271 898
rect 9305 864 9313 898
rect 9263 739 9313 864
rect 9349 1411 9357 1445
rect 9391 1411 9399 1445
rect 9349 1034 9399 1411
rect 9349 1000 9357 1034
rect 9391 1000 9399 1034
rect 9349 966 9399 1000
rect 9349 932 9357 966
rect 9391 932 9399 966
rect 9349 898 9399 932
rect 9349 864 9357 898
rect 9391 864 9399 898
rect 9349 739 9399 864
rect 9435 1361 9485 1445
rect 9435 1327 9443 1361
rect 9477 1327 9485 1361
rect 9435 1034 9485 1327
rect 9435 1000 9443 1034
rect 9477 1000 9485 1034
rect 9435 966 9485 1000
rect 9435 932 9443 966
rect 9477 932 9485 966
rect 9435 898 9485 932
rect 9435 864 9443 898
rect 9477 864 9485 898
rect 9435 739 9485 864
rect 9521 1411 9529 1445
rect 9563 1411 9571 1445
rect 9521 1034 9571 1411
rect 9521 1000 9529 1034
rect 9563 1000 9571 1034
rect 9521 966 9571 1000
rect 9521 932 9529 966
rect 9563 932 9571 966
rect 9521 898 9571 932
rect 9521 864 9529 898
rect 9563 864 9571 898
rect 9521 739 9571 864
rect 9607 1361 9657 1445
rect 9607 1327 9615 1361
rect 9649 1327 9657 1361
rect 9607 1034 9657 1327
rect 9607 1000 9615 1034
rect 9649 1000 9657 1034
rect 9607 966 9657 1000
rect 9607 932 9615 966
rect 9649 932 9657 966
rect 9607 898 9657 932
rect 9607 864 9615 898
rect 9649 864 9657 898
rect 9607 739 9657 864
rect 9693 1411 9701 1445
rect 9735 1411 9743 1445
rect 9693 1034 9743 1411
rect 9693 1000 9701 1034
rect 9735 1000 9743 1034
rect 9693 966 9743 1000
rect 9693 932 9701 966
rect 9735 932 9743 966
rect 9693 898 9743 932
rect 9693 864 9701 898
rect 9735 864 9743 898
rect 9693 739 9743 864
rect 9779 1361 9829 1445
rect 9779 1327 9787 1361
rect 9821 1327 9829 1361
rect 9779 1034 9829 1327
rect 9779 1000 9787 1034
rect 9821 1000 9829 1034
rect 9779 966 9829 1000
rect 9779 932 9787 966
rect 9821 932 9829 966
rect 9779 898 9829 932
rect 9779 864 9787 898
rect 9821 864 9829 898
rect 9779 739 9829 864
rect 9865 1411 9873 1445
rect 9907 1411 9915 1445
rect 9865 1034 9915 1411
rect 9865 1000 9873 1034
rect 9907 1000 9915 1034
rect 9865 966 9915 1000
rect 9865 932 9873 966
rect 9907 932 9915 966
rect 9865 898 9915 932
rect 9865 864 9873 898
rect 9907 864 9915 898
rect 9865 739 9915 864
rect 9951 1361 10001 1445
rect 9951 1327 9959 1361
rect 9993 1327 10001 1361
rect 9951 1034 10001 1327
rect 9951 1000 9959 1034
rect 9993 1000 10001 1034
rect 9951 966 10001 1000
rect 9951 932 9959 966
rect 9993 932 10001 966
rect 9951 898 10001 932
rect 9951 864 9959 898
rect 9993 864 10001 898
rect 9951 739 10001 864
rect 10037 1411 10045 1445
rect 10079 1411 10087 1445
rect 10037 1034 10087 1411
rect 10037 1000 10045 1034
rect 10079 1000 10087 1034
rect 10037 966 10087 1000
rect 10037 932 10045 966
rect 10079 932 10087 966
rect 10037 898 10087 932
rect 10037 864 10045 898
rect 10079 864 10087 898
rect 10037 739 10087 864
rect 10123 1361 10173 1445
rect 10123 1327 10131 1361
rect 10165 1327 10173 1361
rect 10123 1034 10173 1327
rect 10123 1000 10131 1034
rect 10165 1000 10173 1034
rect 10123 966 10173 1000
rect 10123 932 10131 966
rect 10165 932 10173 966
rect 10123 898 10173 932
rect 10123 864 10131 898
rect 10165 864 10173 898
rect 10123 739 10173 864
rect 10209 1411 10217 1445
rect 10251 1411 10259 1445
rect 10209 1034 10259 1411
rect 10209 1000 10217 1034
rect 10251 1000 10259 1034
rect 10209 966 10259 1000
rect 10209 932 10217 966
rect 10251 932 10259 966
rect 10209 898 10259 932
rect 10209 864 10217 898
rect 10251 864 10259 898
rect 10209 739 10259 864
rect 10295 1361 10345 1445
rect 10295 1327 10303 1361
rect 10337 1327 10345 1361
rect 10295 1034 10345 1327
rect 10295 1000 10303 1034
rect 10337 1000 10345 1034
rect 10295 966 10345 1000
rect 10295 932 10303 966
rect 10337 932 10345 966
rect 10295 898 10345 932
rect 10295 864 10303 898
rect 10337 864 10345 898
rect 10295 739 10345 864
rect 10381 1411 10389 1445
rect 10423 1411 10431 1445
rect 10381 1034 10431 1411
rect 10381 1000 10389 1034
rect 10423 1000 10431 1034
rect 10381 966 10431 1000
rect 10381 932 10389 966
rect 10423 932 10431 966
rect 10381 898 10431 932
rect 10381 864 10389 898
rect 10423 864 10431 898
rect 10381 739 10431 864
rect 10467 1361 10517 1445
rect 10467 1327 10475 1361
rect 10509 1327 10517 1361
rect 10467 1034 10517 1327
rect 10467 1000 10475 1034
rect 10509 1000 10517 1034
rect 10467 966 10517 1000
rect 10467 932 10475 966
rect 10509 932 10517 966
rect 10467 898 10517 932
rect 10467 864 10475 898
rect 10509 864 10517 898
rect 10467 739 10517 864
rect 10553 1411 10561 1445
rect 10595 1411 10603 1445
rect 10553 1034 10603 1411
rect 10553 1000 10561 1034
rect 10595 1000 10603 1034
rect 10553 966 10603 1000
rect 10553 932 10561 966
rect 10595 932 10603 966
rect 10553 898 10603 932
rect 10553 864 10561 898
rect 10595 864 10603 898
rect 10553 739 10603 864
rect 10639 1361 10689 1445
rect 10639 1327 10647 1361
rect 10681 1327 10689 1361
rect 10639 1034 10689 1327
rect 10639 1000 10647 1034
rect 10681 1000 10689 1034
rect 10639 966 10689 1000
rect 10639 932 10647 966
rect 10681 932 10689 966
rect 10639 898 10689 932
rect 10639 864 10647 898
rect 10681 864 10689 898
rect 10639 739 10689 864
rect 10725 1411 10733 1445
rect 10767 1411 10775 1445
rect 10725 1034 10775 1411
rect 10725 1000 10733 1034
rect 10767 1000 10775 1034
rect 10725 966 10775 1000
rect 10725 932 10733 966
rect 10767 932 10775 966
rect 10725 898 10775 932
rect 10725 864 10733 898
rect 10767 864 10775 898
rect 10725 739 10775 864
rect 10811 1361 10861 1445
rect 10811 1327 10819 1361
rect 10853 1327 10861 1361
rect 10811 1034 10861 1327
rect 10811 1000 10819 1034
rect 10853 1000 10861 1034
rect 10811 966 10861 1000
rect 10811 932 10819 966
rect 10853 932 10861 966
rect 10811 898 10861 932
rect 10811 864 10819 898
rect 10853 864 10861 898
rect 10811 739 10861 864
rect 10897 1411 10905 1445
rect 10939 1411 10947 1445
rect 10897 1034 10947 1411
rect 10897 1000 10905 1034
rect 10939 1000 10947 1034
rect 10897 966 10947 1000
rect 10897 932 10905 966
rect 10939 932 10947 966
rect 10897 898 10947 932
rect 10897 864 10905 898
rect 10939 864 10947 898
rect 10897 739 10947 864
rect 10983 1361 11033 1445
rect 10983 1327 10991 1361
rect 11025 1327 11033 1361
rect 10983 1034 11033 1327
rect 10983 1000 10991 1034
rect 11025 1000 11033 1034
rect 10983 966 11033 1000
rect 10983 932 10991 966
rect 11025 932 11033 966
rect 10983 898 11033 932
rect 10983 864 10991 898
rect 11025 864 11033 898
rect 10983 739 11033 864
rect 11069 1411 11077 1445
rect 11111 1411 11119 1445
rect 11069 1034 11119 1411
rect 11069 1000 11077 1034
rect 11111 1000 11119 1034
rect 11069 966 11119 1000
rect 11069 932 11077 966
rect 11111 932 11119 966
rect 11069 898 11119 932
rect 11069 864 11077 898
rect 11111 864 11119 898
rect 11069 739 11119 864
rect 11155 1361 11205 1445
rect 11155 1327 11163 1361
rect 11197 1327 11205 1361
rect 11155 1034 11205 1327
rect 11155 1000 11163 1034
rect 11197 1000 11205 1034
rect 11155 966 11205 1000
rect 11155 932 11163 966
rect 11197 932 11205 966
rect 11155 898 11205 932
rect 11155 864 11163 898
rect 11197 864 11205 898
rect 11155 739 11205 864
rect 11241 1411 11249 1445
rect 11283 1411 11291 1445
rect 11241 1034 11291 1411
rect 11241 1000 11249 1034
rect 11283 1000 11291 1034
rect 11241 966 11291 1000
rect 11241 932 11249 966
rect 11283 932 11291 966
rect 11241 898 11291 932
rect 11241 864 11249 898
rect 11283 864 11291 898
rect 11241 739 11291 864
rect 11327 1361 11377 1445
rect 11327 1327 11335 1361
rect 11369 1327 11377 1361
rect 11327 1034 11377 1327
rect 11327 1000 11335 1034
rect 11369 1000 11377 1034
rect 11327 966 11377 1000
rect 11327 932 11335 966
rect 11369 932 11377 966
rect 11327 898 11377 932
rect 11327 864 11335 898
rect 11369 864 11377 898
rect 11327 739 11377 864
rect 233 605 283 689
rect 233 571 241 605
rect 275 571 283 605
rect 233 487 283 571
rect 405 605 455 689
rect 405 571 413 605
rect 447 571 455 605
rect 405 487 455 571
rect 577 605 627 689
rect 577 571 585 605
rect 619 571 627 605
rect 577 487 627 571
rect 749 605 799 689
rect 749 571 757 605
rect 791 571 799 605
rect 749 487 799 571
rect 921 605 971 689
rect 921 571 929 605
rect 963 571 971 605
rect 921 487 971 571
rect 1093 605 1143 689
rect 1093 571 1101 605
rect 1135 571 1143 605
rect 1093 487 1143 571
rect 1265 605 1315 689
rect 1265 571 1273 605
rect 1307 571 1315 605
rect 1265 487 1315 571
rect 1437 605 1487 689
rect 1437 571 1445 605
rect 1479 571 1487 605
rect 1437 487 1487 571
rect 1609 605 1659 689
rect 1609 571 1617 605
rect 1651 571 1659 605
rect 1609 487 1659 571
rect 1781 605 1831 689
rect 1781 571 1789 605
rect 1823 571 1831 605
rect 1781 487 1831 571
rect 1953 605 2003 689
rect 1953 571 1961 605
rect 1995 571 2003 605
rect 1953 487 2003 571
rect 2125 605 2175 689
rect 2125 571 2133 605
rect 2167 571 2175 605
rect 2125 487 2175 571
rect 2641 605 2691 689
rect 2641 571 2649 605
rect 2683 571 2691 605
rect 2641 487 2691 571
rect 2813 605 2863 689
rect 2813 571 2821 605
rect 2855 571 2863 605
rect 2813 487 2863 571
rect 2985 605 3035 689
rect 2985 571 2993 605
rect 3027 571 3035 605
rect 2985 487 3035 571
rect 3157 605 3207 689
rect 3157 571 3165 605
rect 3199 571 3207 605
rect 3157 487 3207 571
rect 3329 605 3379 689
rect 3329 571 3337 605
rect 3371 571 3379 605
rect 3329 487 3379 571
rect 3501 605 3551 689
rect 3501 571 3509 605
rect 3543 571 3551 605
rect 3501 487 3551 571
rect 4017 605 4067 689
rect 4017 571 4025 605
rect 4059 571 4067 605
rect 4017 487 4067 571
rect 4189 605 4239 689
rect 4189 571 4197 605
rect 4231 571 4239 605
rect 4189 487 4239 571
rect 4361 605 4411 689
rect 4361 571 4369 605
rect 4403 571 4411 605
rect 4361 487 4411 571
rect 4533 605 4583 689
rect 4533 571 4541 605
rect 4575 571 4583 605
rect 4533 487 4583 571
rect 4705 605 4755 689
rect 4705 571 4713 605
rect 4747 571 4755 605
rect 4705 487 4755 571
rect 4877 605 4927 689
rect 4877 571 4885 605
rect 4919 571 4927 605
rect 4877 487 4927 571
rect 5393 605 5443 689
rect 5393 571 5401 605
rect 5435 571 5443 605
rect 5393 487 5443 571
rect 5565 605 5615 689
rect 5565 571 5573 605
rect 5607 571 5615 605
rect 5565 487 5615 571
rect 5737 605 5787 689
rect 5737 571 5745 605
rect 5779 571 5787 605
rect 5737 487 5787 571
rect 7285 605 7335 689
rect 7285 571 7293 605
rect 7327 571 7335 605
rect 7285 487 7335 571
rect 7457 605 7507 689
rect 7457 571 7465 605
rect 7499 571 7507 605
rect 7457 487 7507 571
rect 7629 605 7679 689
rect 7629 571 7637 605
rect 7671 571 7679 605
rect 7629 487 7679 571
rect 7801 605 7851 689
rect 7801 571 7809 605
rect 7843 571 7851 605
rect 7801 487 7851 571
rect 7973 605 8023 689
rect 7973 571 7981 605
rect 8015 571 8023 605
rect 7973 487 8023 571
rect 8145 605 8195 689
rect 8145 571 8153 605
rect 8187 571 8195 605
rect 8145 487 8195 571
rect 8317 605 8367 689
rect 8317 571 8325 605
rect 8359 571 8367 605
rect 8317 487 8367 571
rect 8489 605 8539 689
rect 8489 571 8497 605
rect 8531 571 8539 605
rect 8489 487 8539 571
rect 8661 605 8711 689
rect 8661 571 8669 605
rect 8703 571 8711 605
rect 8661 487 8711 571
rect 8833 605 8883 689
rect 8833 571 8841 605
rect 8875 571 8883 605
rect 8833 487 8883 571
rect 9005 605 9055 689
rect 9005 571 9013 605
rect 9047 571 9055 605
rect 9005 487 9055 571
rect 9177 605 9227 689
rect 9177 571 9185 605
rect 9219 571 9227 605
rect 9177 487 9227 571
rect 9349 605 9399 689
rect 9349 571 9357 605
rect 9391 571 9399 605
rect 9349 487 9399 571
rect 9521 605 9571 689
rect 9521 571 9529 605
rect 9563 571 9571 605
rect 9521 487 9571 571
rect 9693 605 9743 689
rect 9693 571 9701 605
rect 9735 571 9743 605
rect 9693 487 9743 571
rect 9865 605 9915 689
rect 9865 571 9873 605
rect 9907 571 9915 605
rect 9865 487 9915 571
rect 10037 605 10087 689
rect 10037 571 10045 605
rect 10079 571 10087 605
rect 10037 487 10087 571
rect 10209 605 10259 689
rect 10209 571 10217 605
rect 10251 571 10259 605
rect 10209 487 10259 571
rect 10381 605 10431 689
rect 10381 571 10389 605
rect 10423 571 10431 605
rect 10381 487 10431 571
rect 10553 605 10603 689
rect 10553 571 10561 605
rect 10595 571 10603 605
rect 10553 487 10603 571
rect 10725 605 10775 689
rect 10725 571 10733 605
rect 10767 571 10775 605
rect 10725 487 10775 571
rect 10897 605 10947 689
rect 10897 571 10905 605
rect 10939 571 10947 605
rect 10897 487 10947 571
rect 11069 605 11119 689
rect 11069 571 11077 605
rect 11111 571 11119 605
rect 11069 487 11119 571
rect 11241 605 11291 689
rect 11241 571 11249 605
rect 11283 571 11291 605
rect 11241 487 11291 571
rect 233 185 283 269
rect 233 151 241 185
rect 275 151 283 185
rect 233 67 283 151
rect 405 185 455 269
rect 405 151 413 185
rect 447 151 455 185
rect 405 67 455 151
rect 577 185 627 269
rect 577 151 585 185
rect 619 151 627 185
rect 577 67 627 151
rect 749 185 799 269
rect 749 151 757 185
rect 791 151 799 185
rect 749 67 799 151
rect 921 185 971 269
rect 921 151 929 185
rect 963 151 971 185
rect 921 67 971 151
rect 1093 185 1143 269
rect 1093 151 1101 185
rect 1135 151 1143 185
rect 1093 67 1143 151
rect 1265 185 1315 269
rect 1265 151 1273 185
rect 1307 151 1315 185
rect 1265 67 1315 151
rect 1437 185 1487 269
rect 1437 151 1445 185
rect 1479 151 1487 185
rect 1437 67 1487 151
rect 1609 185 1659 269
rect 1609 151 1617 185
rect 1651 151 1659 185
rect 1609 67 1659 151
rect 1781 185 1831 269
rect 1781 151 1789 185
rect 1823 151 1831 185
rect 1781 67 1831 151
rect 1953 185 2003 269
rect 1953 151 1961 185
rect 1995 151 2003 185
rect 1953 67 2003 151
rect 2125 185 2175 269
rect 2125 151 2133 185
rect 2167 151 2175 185
rect 2125 67 2175 151
rect 2641 185 2691 269
rect 2641 151 2649 185
rect 2683 151 2691 185
rect 2641 67 2691 151
rect 2813 185 2863 269
rect 2813 151 2821 185
rect 2855 151 2863 185
rect 2813 67 2863 151
rect 2985 185 3035 269
rect 2985 151 2993 185
rect 3027 151 3035 185
rect 2985 67 3035 151
rect 3157 185 3207 269
rect 3157 151 3165 185
rect 3199 151 3207 185
rect 3157 67 3207 151
rect 3329 185 3379 269
rect 3329 151 3337 185
rect 3371 151 3379 185
rect 3329 67 3379 151
rect 3501 185 3551 269
rect 3501 151 3509 185
rect 3543 151 3551 185
rect 3501 67 3551 151
rect 7285 185 7335 269
rect 7285 151 7293 185
rect 7327 151 7335 185
rect 7285 67 7335 151
rect 7457 185 7507 269
rect 7457 151 7465 185
rect 7499 151 7507 185
rect 7457 67 7507 151
rect 7629 185 7679 269
rect 7629 151 7637 185
rect 7671 151 7679 185
rect 7629 67 7679 151
rect 7801 185 7851 269
rect 7801 151 7809 185
rect 7843 151 7851 185
rect 7801 67 7851 151
rect 7973 185 8023 269
rect 7973 151 7981 185
rect 8015 151 8023 185
rect 7973 67 8023 151
rect 8145 185 8195 269
rect 8145 151 8153 185
rect 8187 151 8195 185
rect 8145 67 8195 151
rect 8317 185 8367 269
rect 8317 151 8325 185
rect 8359 151 8367 185
rect 8317 67 8367 151
rect 8489 185 8539 269
rect 8489 151 8497 185
rect 8531 151 8539 185
rect 8489 67 8539 151
rect 8661 185 8711 269
rect 8661 151 8669 185
rect 8703 151 8711 185
rect 8661 67 8711 151
rect 8833 185 8883 269
rect 8833 151 8841 185
rect 8875 151 8883 185
rect 8833 67 8883 151
rect 9005 185 9055 269
rect 9005 151 9013 185
rect 9047 151 9055 185
rect 9005 67 9055 151
rect 9177 185 9227 269
rect 9177 151 9185 185
rect 9219 151 9227 185
rect 9177 67 9227 151
rect 9349 185 9399 269
rect 9349 151 9357 185
rect 9391 151 9399 185
rect 9349 67 9399 151
rect 9521 185 9571 269
rect 9521 151 9529 185
rect 9563 151 9571 185
rect 9521 67 9571 151
rect 9693 185 9743 269
rect 9693 151 9701 185
rect 9735 151 9743 185
rect 9693 67 9743 151
rect 9865 185 9915 269
rect 9865 151 9873 185
rect 9907 151 9915 185
rect 9865 67 9915 151
rect 10037 185 10087 269
rect 10037 151 10045 185
rect 10079 151 10087 185
rect 10037 67 10087 151
rect 10209 185 10259 269
rect 10209 151 10217 185
rect 10251 151 10259 185
rect 10209 67 10259 151
rect 10381 185 10431 269
rect 10381 151 10389 185
rect 10423 151 10431 185
rect 10381 67 10431 151
rect 10553 185 10603 269
rect 10553 151 10561 185
rect 10595 151 10603 185
rect 10553 67 10603 151
rect 10725 185 10775 269
rect 10725 151 10733 185
rect 10767 151 10775 185
rect 10725 67 10775 151
rect 10897 185 10947 269
rect 10897 151 10905 185
rect 10939 151 10947 185
rect 10897 67 10947 151
rect 11069 185 11119 269
rect 11069 151 11077 185
rect 11111 151 11119 185
rect 11069 67 11119 151
rect 11241 185 11291 269
rect 11241 151 11249 185
rect 11283 151 11291 185
rect 11241 67 11291 151
<< viali >>
rect 1187 4015 1221 4049
rect 3079 4015 3113 4049
rect 6777 4015 6811 4049
rect 9271 4015 9305 4049
rect 1187 3595 1221 3629
rect 3079 3595 3113 3629
rect 6261 3679 6295 3713
rect 6777 3595 6811 3629
rect 9271 3595 9305 3629
rect 1101 2839 1135 2873
rect 1187 2755 1221 2789
rect 1273 2839 1307 2873
rect 2993 2839 3027 2873
rect 3079 2755 3113 2789
rect 4455 3259 4489 3293
rect 5573 3259 5607 3293
rect 6261 3259 6295 3293
rect 6605 3259 6639 3293
rect 3165 2839 3199 2873
rect 4455 2839 4489 2873
rect 5573 2839 5607 2873
rect 155 2503 189 2537
rect 241 2587 275 2621
rect 327 2503 361 2537
rect 413 2587 447 2621
rect 499 2503 533 2537
rect 585 2587 619 2621
rect 671 2503 705 2537
rect 757 2587 791 2621
rect 843 2503 877 2537
rect 929 2587 963 2621
rect 1015 2503 1049 2537
rect 1101 2587 1135 2621
rect 1187 2503 1221 2537
rect 1273 2587 1307 2621
rect 1359 2503 1393 2537
rect 1445 2587 1479 2621
rect 1531 2503 1565 2537
rect 1617 2587 1651 2621
rect 1703 2503 1737 2537
rect 1789 2587 1823 2621
rect 1875 2503 1909 2537
rect 1961 2587 1995 2621
rect 2047 2503 2081 2537
rect 2133 2587 2167 2621
rect 2219 2503 2253 2537
rect 2563 2503 2597 2537
rect 2649 2587 2683 2621
rect 2735 2503 2769 2537
rect 2821 2587 2855 2621
rect 2907 2503 2941 2537
rect 2993 2587 3027 2621
rect 3079 2503 3113 2537
rect 3165 2587 3199 2621
rect 3251 2503 3285 2537
rect 3337 2587 3371 2621
rect 3423 2503 3457 2537
rect 3509 2587 3543 2621
rect 3595 2503 3629 2537
rect 4369 2083 4403 2117
rect 4455 1999 4489 2033
rect 4541 2083 4575 2117
rect 5487 2083 5521 2117
rect 5573 1999 5607 2033
rect 6175 2503 6209 2537
rect 6261 2419 6295 2453
rect 6605 2755 6639 2789
rect 6691 2839 6725 2873
rect 6777 2755 6811 2789
rect 6863 2839 6897 2873
rect 9185 2839 9219 2873
rect 9271 2755 9305 2789
rect 9357 2839 9391 2873
rect 6605 2587 6639 2621
rect 6347 2503 6381 2537
rect 6691 2503 6725 2537
rect 5659 2083 5693 2117
rect 6261 2167 6295 2201
rect 5229 1915 5263 1949
rect 6777 2587 6811 2621
rect 6863 2503 6897 2537
rect 7207 2503 7241 2537
rect 7293 2587 7327 2621
rect 7379 2503 7413 2537
rect 7465 2587 7499 2621
rect 7551 2503 7585 2537
rect 7637 2587 7671 2621
rect 7723 2503 7757 2537
rect 7809 2587 7843 2621
rect 7895 2503 7929 2537
rect 7981 2587 8015 2621
rect 8067 2503 8101 2537
rect 8153 2587 8187 2621
rect 8239 2503 8273 2537
rect 8325 2587 8359 2621
rect 8411 2503 8445 2537
rect 8497 2587 8531 2621
rect 8583 2503 8617 2537
rect 8669 2587 8703 2621
rect 8755 2503 8789 2537
rect 8841 2587 8875 2621
rect 8927 2503 8961 2537
rect 9013 2587 9047 2621
rect 9099 2503 9133 2537
rect 9185 2587 9219 2621
rect 9271 2503 9305 2537
rect 9357 2587 9391 2621
rect 9443 2503 9477 2537
rect 9529 2587 9563 2621
rect 9615 2503 9649 2537
rect 9701 2587 9735 2621
rect 9787 2503 9821 2537
rect 9873 2587 9907 2621
rect 9959 2503 9993 2537
rect 10045 2587 10079 2621
rect 10131 2503 10165 2537
rect 10217 2587 10251 2621
rect 10303 2503 10337 2537
rect 10389 2587 10423 2621
rect 10475 2503 10509 2537
rect 10561 2587 10595 2621
rect 10647 2503 10681 2537
rect 10733 2587 10767 2621
rect 10819 2503 10853 2537
rect 10905 2587 10939 2621
rect 10991 2503 11025 2537
rect 11077 2587 11111 2621
rect 11163 2503 11197 2537
rect 11249 2587 11283 2621
rect 11335 2503 11369 2537
rect 241 1747 275 1781
rect 413 1747 447 1781
rect 585 1747 619 1781
rect 757 1747 791 1781
rect 929 1747 963 1781
rect 1101 1747 1135 1781
rect 1273 1747 1307 1781
rect 1445 1747 1479 1781
rect 1617 1747 1651 1781
rect 1789 1747 1823 1781
rect 1961 1747 1995 1781
rect 2133 1747 2167 1781
rect 2649 1747 2683 1781
rect 2821 1747 2855 1781
rect 2993 1747 3027 1781
rect 3165 1747 3199 1781
rect 3337 1747 3371 1781
rect 3509 1747 3543 1781
rect 3939 1747 3973 1781
rect 155 1327 189 1361
rect 241 1411 275 1445
rect 327 1327 361 1361
rect 413 1411 447 1445
rect 499 1327 533 1361
rect 585 1411 619 1445
rect 671 1327 705 1361
rect 757 1411 791 1445
rect 843 1327 877 1361
rect 929 1411 963 1445
rect 1015 1327 1049 1361
rect 1101 1411 1135 1445
rect 1187 1327 1221 1361
rect 1273 1411 1307 1445
rect 1359 1327 1393 1361
rect 1445 1411 1479 1445
rect 1531 1327 1565 1361
rect 1617 1411 1651 1445
rect 1703 1327 1737 1361
rect 1789 1411 1823 1445
rect 1875 1327 1909 1361
rect 1961 1411 1995 1445
rect 2047 1327 2081 1361
rect 2133 1411 2167 1445
rect 2219 1327 2253 1361
rect 2563 1327 2597 1361
rect 2649 1411 2683 1445
rect 2735 1327 2769 1361
rect 2821 1411 2855 1445
rect 2907 1327 2941 1361
rect 2993 1411 3027 1445
rect 3079 1327 3113 1361
rect 3165 1411 3199 1445
rect 3251 1327 3285 1361
rect 3337 1411 3371 1445
rect 3423 1327 3457 1361
rect 3509 1411 3543 1445
rect 3595 1327 3629 1361
rect 4025 1831 4059 1865
rect 4111 1747 4145 1781
rect 4197 1831 4231 1865
rect 4283 1747 4317 1781
rect 4369 1831 4403 1865
rect 4455 1747 4489 1781
rect 4541 1831 4575 1865
rect 4627 1747 4661 1781
rect 4713 1831 4747 1865
rect 4799 1747 4833 1781
rect 4885 1831 4919 1865
rect 5229 1831 5263 1865
rect 4971 1747 5005 1781
rect 5315 1747 5349 1781
rect 5401 1831 5435 1865
rect 5487 1747 5521 1781
rect 5573 1831 5607 1865
rect 5659 1747 5693 1781
rect 5745 1831 5779 1865
rect 5831 1747 5865 1781
rect 6261 1747 6295 1781
rect 6777 1747 6811 1781
rect 7293 1747 7327 1781
rect 7465 1747 7499 1781
rect 7637 1747 7671 1781
rect 7809 1747 7843 1781
rect 7981 1747 8015 1781
rect 8153 1747 8187 1781
rect 8325 1747 8359 1781
rect 8497 1747 8531 1781
rect 8669 1747 8703 1781
rect 8841 1747 8875 1781
rect 9013 1747 9047 1781
rect 9185 1747 9219 1781
rect 9357 1747 9391 1781
rect 9529 1747 9563 1781
rect 9701 1747 9735 1781
rect 9873 1747 9907 1781
rect 10045 1747 10079 1781
rect 10217 1747 10251 1781
rect 10389 1747 10423 1781
rect 10561 1747 10595 1781
rect 10733 1747 10767 1781
rect 10905 1747 10939 1781
rect 11077 1747 11111 1781
rect 11249 1747 11283 1781
rect 4025 991 4059 1025
rect 4197 991 4231 1025
rect 4369 991 4403 1025
rect 4541 991 4575 1025
rect 4713 991 4747 1025
rect 4885 991 4919 1025
rect 5401 991 5435 1025
rect 5573 991 5607 1025
rect 5745 991 5779 1025
rect 6175 991 6209 1025
rect 6261 907 6295 941
rect 6777 1327 6811 1361
rect 7207 1327 7241 1361
rect 6347 991 6381 1025
rect 7293 1411 7327 1445
rect 7379 1327 7413 1361
rect 7465 1411 7499 1445
rect 7551 1327 7585 1361
rect 7637 1411 7671 1445
rect 7723 1327 7757 1361
rect 7809 1411 7843 1445
rect 7895 1327 7929 1361
rect 7981 1411 8015 1445
rect 8067 1327 8101 1361
rect 8153 1411 8187 1445
rect 8239 1327 8273 1361
rect 8325 1411 8359 1445
rect 8411 1327 8445 1361
rect 8497 1411 8531 1445
rect 8583 1327 8617 1361
rect 8669 1411 8703 1445
rect 8755 1327 8789 1361
rect 8841 1411 8875 1445
rect 8927 1327 8961 1361
rect 9013 1411 9047 1445
rect 9099 1327 9133 1361
rect 9185 1411 9219 1445
rect 9271 1327 9305 1361
rect 9357 1411 9391 1445
rect 9443 1327 9477 1361
rect 9529 1411 9563 1445
rect 9615 1327 9649 1361
rect 9701 1411 9735 1445
rect 9787 1327 9821 1361
rect 9873 1411 9907 1445
rect 9959 1327 9993 1361
rect 10045 1411 10079 1445
rect 10131 1327 10165 1361
rect 10217 1411 10251 1445
rect 10303 1327 10337 1361
rect 10389 1411 10423 1445
rect 10475 1327 10509 1361
rect 10561 1411 10595 1445
rect 10647 1327 10681 1361
rect 10733 1411 10767 1445
rect 10819 1327 10853 1361
rect 10905 1411 10939 1445
rect 10991 1327 11025 1361
rect 11077 1411 11111 1445
rect 11163 1327 11197 1361
rect 11249 1411 11283 1445
rect 11335 1327 11369 1361
rect 241 571 275 605
rect 413 571 447 605
rect 585 571 619 605
rect 757 571 791 605
rect 929 571 963 605
rect 1101 571 1135 605
rect 1273 571 1307 605
rect 1445 571 1479 605
rect 1617 571 1651 605
rect 1789 571 1823 605
rect 1961 571 1995 605
rect 2133 571 2167 605
rect 2649 571 2683 605
rect 2821 571 2855 605
rect 2993 571 3027 605
rect 3165 571 3199 605
rect 3337 571 3371 605
rect 3509 571 3543 605
rect 4025 571 4059 605
rect 4197 571 4231 605
rect 4369 571 4403 605
rect 4541 571 4575 605
rect 4713 571 4747 605
rect 4885 571 4919 605
rect 5401 571 5435 605
rect 5573 571 5607 605
rect 5745 571 5779 605
rect 7293 571 7327 605
rect 7465 571 7499 605
rect 7637 571 7671 605
rect 7809 571 7843 605
rect 7981 571 8015 605
rect 8153 571 8187 605
rect 8325 571 8359 605
rect 8497 571 8531 605
rect 8669 571 8703 605
rect 8841 571 8875 605
rect 9013 571 9047 605
rect 9185 571 9219 605
rect 9357 571 9391 605
rect 9529 571 9563 605
rect 9701 571 9735 605
rect 9873 571 9907 605
rect 10045 571 10079 605
rect 10217 571 10251 605
rect 10389 571 10423 605
rect 10561 571 10595 605
rect 10733 571 10767 605
rect 10905 571 10939 605
rect 11077 571 11111 605
rect 11249 571 11283 605
rect 241 151 275 185
rect 413 151 447 185
rect 585 151 619 185
rect 757 151 791 185
rect 929 151 963 185
rect 1101 151 1135 185
rect 1273 151 1307 185
rect 1445 151 1479 185
rect 1617 151 1651 185
rect 1789 151 1823 185
rect 1961 151 1995 185
rect 2133 151 2167 185
rect 2649 151 2683 185
rect 2821 151 2855 185
rect 2993 151 3027 185
rect 3165 151 3199 185
rect 3337 151 3371 185
rect 3509 151 3543 185
rect 7293 151 7327 185
rect 7465 151 7499 185
rect 7637 151 7671 185
rect 7809 151 7843 185
rect 7981 151 8015 185
rect 8153 151 8187 185
rect 8325 151 8359 185
rect 8497 151 8531 185
rect 8669 151 8703 185
rect 8841 151 8875 185
rect 9013 151 9047 185
rect 9185 151 9219 185
rect 9357 151 9391 185
rect 9529 151 9563 185
rect 9701 151 9735 185
rect 9873 151 9907 185
rect 10045 151 10079 185
rect 10217 151 10251 185
rect 10389 151 10423 185
rect 10561 151 10595 185
rect 10733 151 10767 185
rect 10905 151 10939 185
rect 11077 151 11111 185
rect 11249 151 11283 185
<< metal1 >>
rect 1084 4058 1324 4060
rect 1084 4049 1264 4058
rect 1084 4015 1187 4049
rect 1221 4015 1264 4049
rect 1084 4006 1264 4015
rect 1316 4006 1324 4058
rect 1084 4004 1324 4006
rect 2976 4058 3216 4060
rect 2976 4006 2984 4058
rect 3036 4049 3216 4058
rect 3036 4015 3079 4049
rect 3113 4015 3216 4049
rect 3036 4006 3216 4015
rect 2976 4004 3216 4006
rect 6674 4058 6914 4060
rect 6674 4049 6854 4058
rect 6674 4015 6777 4049
rect 6811 4015 6854 4049
rect 6674 4006 6854 4015
rect 6906 4006 6914 4058
rect 6674 4004 6914 4006
rect 9168 4058 9408 4060
rect 9168 4006 9176 4058
rect 9228 4049 9408 4058
rect 9228 4015 9271 4049
rect 9305 4015 9408 4049
rect 9228 4006 9408 4015
rect 9168 4004 9408 4006
rect 5472 3722 9234 3724
rect 5472 3670 5478 3722
rect 5530 3713 6854 3722
rect 5530 3679 6261 3713
rect 6295 3679 6854 3713
rect 5530 3670 6854 3679
rect 6906 3670 9176 3722
rect 9228 3670 9234 3722
rect 5472 3668 9234 3670
rect 998 3638 1238 3640
rect 998 3586 1178 3638
rect 1230 3586 1238 3638
rect 998 3584 1238 3586
rect 3062 3638 3302 3640
rect 3062 3586 3070 3638
rect 3122 3586 3302 3638
rect 3062 3584 3302 3586
rect 6588 3638 6828 3640
rect 6588 3586 6596 3638
rect 6648 3629 6828 3638
rect 6648 3595 6777 3629
rect 6811 3595 6828 3629
rect 6648 3586 6828 3595
rect 6588 3584 6828 3586
rect 9254 3638 9494 3640
rect 9254 3586 9262 3638
rect 9314 3586 9494 3638
rect 9254 3584 9494 3586
rect 4352 3302 4592 3304
rect 4352 3293 4532 3302
rect 4352 3259 4455 3293
rect 4489 3259 4532 3293
rect 4352 3250 4532 3259
rect 4584 3250 4592 3302
rect 4352 3248 4592 3250
rect 5470 3302 5710 3304
rect 5470 3250 5478 3302
rect 5530 3293 5710 3302
rect 5530 3259 5573 3293
rect 5607 3259 5710 3293
rect 5530 3250 5710 3259
rect 5470 3248 5710 3250
rect 6244 3293 6656 3304
rect 6244 3259 6261 3293
rect 6295 3259 6605 3293
rect 6639 3259 6656 3293
rect 6244 3248 6656 3259
rect 1258 2966 4590 2968
rect 1258 2914 1264 2966
rect 1316 2914 2984 2966
rect 3036 2914 4532 2966
rect 4584 2914 4590 2966
rect 1258 2912 4590 2914
rect 1084 2882 1324 2884
rect 1084 2873 1264 2882
rect 1084 2839 1101 2873
rect 1135 2839 1264 2873
rect 1084 2830 1264 2839
rect 1316 2830 1324 2882
rect 1084 2828 1324 2830
rect 2976 2882 3216 2884
rect 2976 2830 2984 2882
rect 3036 2873 3216 2882
rect 3036 2839 3165 2873
rect 3199 2839 3216 2873
rect 3036 2830 3216 2839
rect 2976 2828 3216 2830
rect 4266 2882 4506 2884
rect 4266 2830 4274 2882
rect 4326 2873 4506 2882
rect 4326 2839 4455 2873
rect 4489 2839 4506 2873
rect 4326 2830 4506 2839
rect 4266 2828 4506 2830
rect 5556 2882 5796 2884
rect 5556 2873 5650 2882
rect 5556 2839 5573 2873
rect 5607 2839 5650 2873
rect 5556 2830 5650 2839
rect 5702 2830 5796 2882
rect 5556 2828 5796 2830
rect 6674 2882 6914 2884
rect 6674 2873 6854 2882
rect 6674 2839 6691 2873
rect 6725 2839 6854 2873
rect 6674 2830 6854 2839
rect 6906 2830 6914 2882
rect 6674 2828 6914 2830
rect 9168 2882 9408 2884
rect 9168 2830 9176 2882
rect 9228 2873 9408 2882
rect 9228 2839 9357 2873
rect 9391 2839 9408 2873
rect 9228 2830 9408 2839
rect 9168 2828 9408 2830
rect 998 2798 2956 2800
rect 998 2746 1092 2798
rect 1144 2789 2898 2798
rect 1144 2755 1187 2789
rect 1221 2755 2898 2789
rect 1144 2746 2898 2755
rect 2950 2746 2956 2798
rect 998 2744 2956 2746
rect 3062 2798 3302 2800
rect 3062 2789 3156 2798
rect 3062 2755 3079 2789
rect 3113 2755 3156 2789
rect 3062 2746 3156 2755
rect 3208 2746 3302 2798
rect 3062 2744 3302 2746
rect 6588 2789 6828 2800
rect 6588 2755 6605 2789
rect 6639 2755 6777 2789
rect 6811 2755 6828 2789
rect 6588 2744 6828 2755
rect 9254 2798 9494 2800
rect 9254 2789 9348 2798
rect 9254 2755 9271 2789
rect 9305 2755 9348 2789
rect 9254 2746 9348 2755
rect 9400 2746 9494 2798
rect 9254 2744 9494 2746
rect 224 2630 2184 2632
rect 224 2621 1092 2630
rect 1144 2621 2184 2630
rect 224 2587 241 2621
rect 275 2587 413 2621
rect 447 2587 585 2621
rect 619 2587 757 2621
rect 791 2587 929 2621
rect 963 2587 1092 2621
rect 1144 2587 1273 2621
rect 1307 2587 1445 2621
rect 1479 2587 1617 2621
rect 1651 2587 1789 2621
rect 1823 2587 1961 2621
rect 1995 2587 2133 2621
rect 2167 2587 2184 2621
rect 224 2578 1092 2587
rect 1144 2578 2184 2587
rect 224 2576 2184 2578
rect 2632 2630 3560 2632
rect 2632 2621 3156 2630
rect 3208 2621 3560 2630
rect 2632 2587 2649 2621
rect 2683 2587 2821 2621
rect 2855 2587 2993 2621
rect 3027 2587 3156 2621
rect 3208 2587 3337 2621
rect 3371 2587 3509 2621
rect 3543 2587 3560 2621
rect 2632 2578 3156 2587
rect 3208 2578 3560 2587
rect 2632 2576 3560 2578
rect 6588 2621 6828 2632
rect 6588 2587 6605 2621
rect 6639 2587 6777 2621
rect 6811 2587 6828 2621
rect 6588 2576 6828 2587
rect 7276 2630 11300 2632
rect 7276 2621 9348 2630
rect 9400 2621 11300 2630
rect 7276 2587 7293 2621
rect 7327 2587 7465 2621
rect 7499 2587 7637 2621
rect 7671 2587 7809 2621
rect 7843 2587 7981 2621
rect 8015 2587 8153 2621
rect 8187 2587 8325 2621
rect 8359 2587 8497 2621
rect 8531 2587 8669 2621
rect 8703 2587 8841 2621
rect 8875 2587 9013 2621
rect 9047 2587 9185 2621
rect 9219 2587 9348 2621
rect 9400 2587 9529 2621
rect 9563 2587 9701 2621
rect 9735 2587 9873 2621
rect 9907 2587 10045 2621
rect 10079 2587 10217 2621
rect 10251 2587 10389 2621
rect 10423 2587 10561 2621
rect 10595 2587 10733 2621
rect 10767 2587 10905 2621
rect 10939 2587 11077 2621
rect 11111 2587 11249 2621
rect 11283 2587 11300 2621
rect 7276 2578 9348 2587
rect 9400 2578 11300 2587
rect 7276 2576 11300 2578
rect 138 2546 2270 2548
rect 138 2537 1264 2546
rect 138 2503 155 2537
rect 189 2503 327 2537
rect 361 2503 499 2537
rect 533 2503 671 2537
rect 705 2503 843 2537
rect 877 2503 1015 2537
rect 1049 2503 1187 2537
rect 1221 2503 1264 2537
rect 138 2494 1264 2503
rect 1316 2537 2270 2546
rect 1316 2503 1359 2537
rect 1393 2503 1531 2537
rect 1565 2503 1703 2537
rect 1737 2503 1875 2537
rect 1909 2503 2047 2537
rect 2081 2503 2219 2537
rect 2253 2503 2270 2537
rect 1316 2494 2270 2503
rect 138 2492 2270 2494
rect 2546 2546 3646 2548
rect 2546 2537 2984 2546
rect 2546 2503 2563 2537
rect 2597 2503 2735 2537
rect 2769 2503 2907 2537
rect 2941 2503 2984 2537
rect 2546 2494 2984 2503
rect 3036 2537 3646 2546
rect 3036 2503 3079 2537
rect 3113 2503 3251 2537
rect 3285 2503 3423 2537
rect 3457 2503 3595 2537
rect 3629 2503 3646 2537
rect 3036 2494 3646 2503
rect 2546 2492 3646 2494
rect 5644 2546 6398 2548
rect 5644 2494 5650 2546
rect 5702 2537 6398 2546
rect 5702 2503 6175 2537
rect 6209 2503 6347 2537
rect 6381 2503 6398 2537
rect 5702 2494 6398 2503
rect 5644 2492 6398 2494
rect 6674 2546 6914 2548
rect 6674 2537 6854 2546
rect 6674 2503 6691 2537
rect 6725 2503 6854 2537
rect 6674 2494 6854 2503
rect 6906 2494 6914 2546
rect 6674 2492 6914 2494
rect 7190 2546 11386 2548
rect 7190 2537 9176 2546
rect 7190 2503 7207 2537
rect 7241 2503 7379 2537
rect 7413 2503 7551 2537
rect 7585 2503 7723 2537
rect 7757 2503 7895 2537
rect 7929 2503 8067 2537
rect 8101 2503 8239 2537
rect 8273 2503 8411 2537
rect 8445 2503 8583 2537
rect 8617 2503 8755 2537
rect 8789 2503 8927 2537
rect 8961 2503 9099 2537
rect 9133 2503 9176 2537
rect 7190 2494 9176 2503
rect 9228 2537 11386 2546
rect 9228 2503 9271 2537
rect 9305 2503 9443 2537
rect 9477 2503 9615 2537
rect 9649 2503 9787 2537
rect 9821 2503 9959 2537
rect 9993 2503 10131 2537
rect 10165 2503 10303 2537
rect 10337 2503 10475 2537
rect 10509 2503 10647 2537
rect 10681 2503 10819 2537
rect 10853 2503 10991 2537
rect 11025 2503 11163 2537
rect 11197 2503 11335 2537
rect 11369 2503 11386 2537
rect 9228 2494 11386 2503
rect 7190 2492 11386 2494
rect 6244 2462 9406 2464
rect 6244 2453 9348 2462
rect 6244 2419 6261 2453
rect 6295 2419 9348 2453
rect 6244 2410 9348 2419
rect 9400 2410 9406 2462
rect 6244 2408 9406 2410
rect 4526 2210 6484 2212
rect 4526 2158 4532 2210
rect 4584 2158 5478 2210
rect 5530 2201 6484 2210
rect 5530 2167 6261 2201
rect 6295 2167 6484 2201
rect 5530 2158 6484 2167
rect 4526 2156 6484 2158
rect 4352 2126 4592 2128
rect 4352 2117 4532 2126
rect 4352 2083 4369 2117
rect 4403 2083 4532 2117
rect 4352 2074 4532 2083
rect 4584 2074 4592 2126
rect 4352 2072 4592 2074
rect 5470 2126 5710 2128
rect 5470 2074 5478 2126
rect 5530 2117 5710 2126
rect 5530 2083 5659 2117
rect 5693 2083 5710 2117
rect 5530 2074 5710 2083
rect 5470 2072 5710 2074
rect 4266 2042 4506 2044
rect 4266 1990 4360 2042
rect 4412 2033 4506 2042
rect 4412 1999 4455 2033
rect 4489 1999 4506 2033
rect 4412 1990 4506 1999
rect 4266 1988 4506 1990
rect 5556 2042 5796 2044
rect 5556 1990 5564 2042
rect 5616 1990 5796 2042
rect 5556 1988 5796 1990
rect 4268 1958 5280 1960
rect 4268 1906 4274 1958
rect 4326 1949 5280 1958
rect 4326 1915 5229 1949
rect 5263 1915 5280 1949
rect 4326 1906 5280 1915
rect 4268 1904 5280 1906
rect 3064 1874 4936 1876
rect 3064 1822 3070 1874
rect 3122 1865 4360 1874
rect 4412 1865 4936 1874
rect 3122 1831 4025 1865
rect 4059 1831 4197 1865
rect 4231 1831 4360 1865
rect 4412 1831 4541 1865
rect 4575 1831 4713 1865
rect 4747 1831 4885 1865
rect 4919 1831 4936 1865
rect 3122 1822 4360 1831
rect 4412 1822 4936 1831
rect 3064 1820 4936 1822
rect 5212 1874 5796 1876
rect 5212 1865 5564 1874
rect 5616 1865 5796 1874
rect 5212 1831 5229 1865
rect 5263 1831 5401 1865
rect 5435 1831 5564 1865
rect 5616 1831 5745 1865
rect 5779 1831 5796 1865
rect 5212 1822 5564 1831
rect 5616 1822 5796 1831
rect 5212 1820 5796 1822
rect 224 1790 2184 1792
rect 224 1781 1178 1790
rect 224 1747 241 1781
rect 275 1747 413 1781
rect 447 1747 585 1781
rect 619 1747 757 1781
rect 791 1747 929 1781
rect 963 1747 1101 1781
rect 1135 1747 1178 1781
rect 224 1738 1178 1747
rect 1230 1781 2184 1790
rect 1230 1747 1273 1781
rect 1307 1747 1445 1781
rect 1479 1747 1617 1781
rect 1651 1747 1789 1781
rect 1823 1747 1961 1781
rect 1995 1747 2133 1781
rect 2167 1747 2184 1781
rect 1230 1738 2184 1747
rect 224 1736 2184 1738
rect 2632 1790 3560 1792
rect 2632 1781 3070 1790
rect 2632 1747 2649 1781
rect 2683 1747 2821 1781
rect 2855 1747 2993 1781
rect 3027 1747 3070 1781
rect 2632 1738 3070 1747
rect 3122 1781 3560 1790
rect 3122 1747 3165 1781
rect 3199 1747 3337 1781
rect 3371 1747 3509 1781
rect 3543 1747 3560 1781
rect 3122 1738 3560 1747
rect 2632 1736 3560 1738
rect 3922 1790 5022 1792
rect 3922 1781 4532 1790
rect 3922 1747 3939 1781
rect 3973 1747 4111 1781
rect 4145 1747 4283 1781
rect 4317 1747 4455 1781
rect 4489 1747 4532 1781
rect 3922 1738 4532 1747
rect 4584 1781 5022 1790
rect 4584 1747 4627 1781
rect 4661 1747 4799 1781
rect 4833 1747 4971 1781
rect 5005 1747 5022 1781
rect 4584 1738 5022 1747
rect 3922 1736 5022 1738
rect 5298 1790 5882 1792
rect 5298 1781 5478 1790
rect 5530 1781 5882 1790
rect 5298 1747 5315 1781
rect 5349 1747 5478 1781
rect 5530 1747 5659 1781
rect 5693 1747 5831 1781
rect 5865 1747 5882 1781
rect 5298 1738 5478 1747
rect 5530 1738 5882 1747
rect 5298 1736 5882 1738
rect 6244 1790 6828 1792
rect 6244 1781 6596 1790
rect 6244 1747 6261 1781
rect 6295 1747 6596 1781
rect 6244 1738 6596 1747
rect 6648 1781 6828 1790
rect 6648 1747 6777 1781
rect 6811 1747 6828 1781
rect 6648 1738 6828 1747
rect 6244 1736 6828 1738
rect 7276 1790 11300 1792
rect 7276 1781 9262 1790
rect 7276 1747 7293 1781
rect 7327 1747 7465 1781
rect 7499 1747 7637 1781
rect 7671 1747 7809 1781
rect 7843 1747 7981 1781
rect 8015 1747 8153 1781
rect 8187 1747 8325 1781
rect 8359 1747 8497 1781
rect 8531 1747 8669 1781
rect 8703 1747 8841 1781
rect 8875 1747 9013 1781
rect 9047 1747 9185 1781
rect 9219 1747 9262 1781
rect 7276 1738 9262 1747
rect 9314 1781 11300 1790
rect 9314 1747 9357 1781
rect 9391 1747 9529 1781
rect 9563 1747 9701 1781
rect 9735 1747 9873 1781
rect 9907 1747 10045 1781
rect 10079 1747 10217 1781
rect 10251 1747 10389 1781
rect 10423 1747 10561 1781
rect 10595 1747 10733 1781
rect 10767 1747 10905 1781
rect 10939 1747 11077 1781
rect 11111 1747 11249 1781
rect 11283 1747 11300 1781
rect 9314 1738 11300 1747
rect 7276 1736 11300 1738
rect 1172 1538 3214 1540
rect 1172 1486 1178 1538
rect 1230 1486 3156 1538
rect 3208 1486 3214 1538
rect 1172 1484 3214 1486
rect 224 1454 2184 1456
rect 224 1445 1092 1454
rect 1144 1445 2184 1454
rect 224 1411 241 1445
rect 275 1411 413 1445
rect 447 1411 585 1445
rect 619 1411 757 1445
rect 791 1411 929 1445
rect 963 1411 1092 1445
rect 1144 1411 1273 1445
rect 1307 1411 1445 1445
rect 1479 1411 1617 1445
rect 1651 1411 1789 1445
rect 1823 1411 1961 1445
rect 1995 1411 2133 1445
rect 2167 1411 2184 1445
rect 224 1402 1092 1411
rect 1144 1402 2184 1411
rect 224 1400 2184 1402
rect 2632 1454 3560 1456
rect 2632 1445 3156 1454
rect 3208 1445 3560 1454
rect 2632 1411 2649 1445
rect 2683 1411 2821 1445
rect 2855 1411 2993 1445
rect 3027 1411 3156 1445
rect 3208 1411 3337 1445
rect 3371 1411 3509 1445
rect 3543 1411 3560 1445
rect 2632 1402 3156 1411
rect 3208 1402 3560 1411
rect 2632 1400 3560 1402
rect 7276 1454 11300 1456
rect 7276 1445 9348 1454
rect 9400 1445 11300 1454
rect 7276 1411 7293 1445
rect 7327 1411 7465 1445
rect 7499 1411 7637 1445
rect 7671 1411 7809 1445
rect 7843 1411 7981 1445
rect 8015 1411 8153 1445
rect 8187 1411 8325 1445
rect 8359 1411 8497 1445
rect 8531 1411 8669 1445
rect 8703 1411 8841 1445
rect 8875 1411 9013 1445
rect 9047 1411 9185 1445
rect 9219 1411 9348 1445
rect 9400 1411 9529 1445
rect 9563 1411 9701 1445
rect 9735 1411 9873 1445
rect 9907 1411 10045 1445
rect 10079 1411 10217 1445
rect 10251 1411 10389 1445
rect 10423 1411 10561 1445
rect 10595 1411 10733 1445
rect 10767 1411 10905 1445
rect 10939 1411 11077 1445
rect 11111 1411 11249 1445
rect 11283 1411 11300 1445
rect 7276 1402 9348 1411
rect 9400 1402 11300 1411
rect 7276 1400 11300 1402
rect 138 1370 2270 1372
rect 138 1361 1264 1370
rect 138 1327 155 1361
rect 189 1327 327 1361
rect 361 1327 499 1361
rect 533 1327 671 1361
rect 705 1327 843 1361
rect 877 1327 1015 1361
rect 1049 1327 1187 1361
rect 1221 1327 1264 1361
rect 138 1318 1264 1327
rect 1316 1361 2270 1370
rect 1316 1327 1359 1361
rect 1393 1327 1531 1361
rect 1565 1327 1703 1361
rect 1737 1327 1875 1361
rect 1909 1327 2047 1361
rect 2081 1327 2219 1361
rect 2253 1327 2270 1361
rect 1316 1318 2270 1327
rect 138 1316 2270 1318
rect 2546 1370 3646 1372
rect 2546 1361 2984 1370
rect 2546 1327 2563 1361
rect 2597 1327 2735 1361
rect 2769 1327 2907 1361
rect 2941 1327 2984 1361
rect 2546 1318 2984 1327
rect 3036 1361 3646 1370
rect 3036 1327 3079 1361
rect 3113 1327 3251 1361
rect 3285 1327 3423 1361
rect 3457 1327 3595 1361
rect 3629 1327 3646 1361
rect 3036 1318 3646 1327
rect 2546 1316 3646 1318
rect 6674 1370 6914 1372
rect 6674 1361 6854 1370
rect 6674 1327 6777 1361
rect 6811 1327 6854 1361
rect 6674 1318 6854 1327
rect 6906 1318 6914 1370
rect 6674 1316 6914 1318
rect 7190 1370 11386 1372
rect 7190 1361 9176 1370
rect 7190 1327 7207 1361
rect 7241 1327 7379 1361
rect 7413 1327 7551 1361
rect 7585 1327 7723 1361
rect 7757 1327 7895 1361
rect 7929 1327 8067 1361
rect 8101 1327 8239 1361
rect 8273 1327 8411 1361
rect 8445 1327 8583 1361
rect 8617 1327 8755 1361
rect 8789 1327 8927 1361
rect 8961 1327 9099 1361
rect 9133 1327 9176 1361
rect 7190 1318 9176 1327
rect 9228 1361 11386 1370
rect 9228 1327 9271 1361
rect 9305 1327 9443 1361
rect 9477 1327 9615 1361
rect 9649 1327 9787 1361
rect 9821 1327 9959 1361
rect 9993 1327 10131 1361
rect 10165 1327 10303 1361
rect 10337 1327 10475 1361
rect 10509 1327 10647 1361
rect 10681 1327 10819 1361
rect 10853 1327 10991 1361
rect 11025 1327 11163 1361
rect 11197 1327 11335 1361
rect 11369 1327 11386 1361
rect 9228 1318 11386 1327
rect 7190 1316 11386 1318
rect 4008 1034 4936 1036
rect 4008 1025 4274 1034
rect 4008 991 4025 1025
rect 4059 991 4197 1025
rect 4231 991 4274 1025
rect 4008 982 4274 991
rect 4326 1025 4936 1034
rect 4326 991 4369 1025
rect 4403 991 4541 1025
rect 4575 991 4713 1025
rect 4747 991 4885 1025
rect 4919 991 4936 1025
rect 4326 982 4936 991
rect 4008 980 4936 982
rect 5384 1034 6398 1036
rect 5384 1025 5650 1034
rect 5384 991 5401 1025
rect 5435 991 5573 1025
rect 5607 991 5650 1025
rect 5384 982 5650 991
rect 5702 1025 6398 1034
rect 5702 991 5745 1025
rect 5779 991 6175 1025
rect 6209 991 6347 1025
rect 6381 991 6398 1025
rect 5702 982 6398 991
rect 5384 980 6398 982
rect 5472 950 9234 952
rect 5472 898 5478 950
rect 5530 941 6854 950
rect 5530 907 6261 941
rect 6295 907 6854 941
rect 5530 898 6854 907
rect 6906 898 9176 950
rect 9228 898 9234 950
rect 5472 896 9234 898
rect 2978 698 5536 700
rect 2978 646 2984 698
rect 3036 646 4532 698
rect 4584 646 5478 698
rect 5530 646 5536 698
rect 2978 644 5536 646
rect 224 614 2184 616
rect 224 605 1178 614
rect 224 571 241 605
rect 275 571 413 605
rect 447 571 585 605
rect 619 571 757 605
rect 791 571 929 605
rect 963 571 1101 605
rect 1135 571 1178 605
rect 224 562 1178 571
rect 1230 605 2184 614
rect 1230 571 1273 605
rect 1307 571 1445 605
rect 1479 571 1617 605
rect 1651 571 1789 605
rect 1823 571 1961 605
rect 1995 571 2133 605
rect 2167 571 2184 605
rect 1230 562 2184 571
rect 224 560 2184 562
rect 2632 614 3560 616
rect 2632 605 3070 614
rect 2632 571 2649 605
rect 2683 571 2821 605
rect 2855 571 2993 605
rect 3027 571 3070 605
rect 2632 562 3070 571
rect 3122 605 3560 614
rect 3122 571 3165 605
rect 3199 571 3337 605
rect 3371 571 3509 605
rect 3543 571 3560 605
rect 3122 562 3560 571
rect 2632 560 3560 562
rect 4008 614 4936 616
rect 4008 605 4532 614
rect 4584 605 4936 614
rect 4008 571 4025 605
rect 4059 571 4197 605
rect 4231 571 4369 605
rect 4403 571 4532 605
rect 4584 571 4713 605
rect 4747 571 4885 605
rect 4919 571 4936 605
rect 4008 562 4532 571
rect 4584 562 4936 571
rect 4008 560 4936 562
rect 5384 614 5796 616
rect 5384 605 5478 614
rect 5384 571 5401 605
rect 5435 571 5478 605
rect 5384 562 5478 571
rect 5530 605 5796 614
rect 5530 571 5573 605
rect 5607 571 5745 605
rect 5779 571 5796 605
rect 5530 562 5796 571
rect 5384 560 5796 562
rect 7276 614 11300 616
rect 7276 605 9262 614
rect 7276 571 7293 605
rect 7327 571 7465 605
rect 7499 571 7637 605
rect 7671 571 7809 605
rect 7843 571 7981 605
rect 8015 571 8153 605
rect 8187 571 8325 605
rect 8359 571 8497 605
rect 8531 571 8669 605
rect 8703 571 8841 605
rect 8875 571 9013 605
rect 9047 571 9185 605
rect 9219 571 9262 605
rect 7276 562 9262 571
rect 9314 605 11300 614
rect 9314 571 9357 605
rect 9391 571 9529 605
rect 9563 571 9701 605
rect 9735 571 9873 605
rect 9907 571 10045 605
rect 10079 571 10217 605
rect 10251 571 10389 605
rect 10423 571 10561 605
rect 10595 571 10733 605
rect 10767 571 10905 605
rect 10939 571 11077 605
rect 11111 571 11249 605
rect 11283 571 11300 605
rect 9314 562 11300 571
rect 7276 560 11300 562
rect 1258 278 3042 280
rect 1258 226 1264 278
rect 1316 226 2984 278
rect 3036 226 3042 278
rect 1258 224 3042 226
rect 224 194 2184 196
rect 224 185 1264 194
rect 1316 185 2184 194
rect 224 151 241 185
rect 275 151 413 185
rect 447 151 585 185
rect 619 151 757 185
rect 791 151 929 185
rect 963 151 1101 185
rect 1135 151 1264 185
rect 1316 151 1445 185
rect 1479 151 1617 185
rect 1651 151 1789 185
rect 1823 151 1961 185
rect 1995 151 2133 185
rect 2167 151 2184 185
rect 224 142 1264 151
rect 1316 142 2184 151
rect 224 140 2184 142
rect 2632 194 3560 196
rect 2632 185 2984 194
rect 3036 185 3560 194
rect 2632 151 2649 185
rect 2683 151 2821 185
rect 2855 151 2984 185
rect 3036 151 3165 185
rect 3199 151 3337 185
rect 3371 151 3509 185
rect 3543 151 3560 185
rect 2632 142 2984 151
rect 3036 142 3560 151
rect 2632 140 3560 142
rect 7276 194 11300 196
rect 7276 185 9176 194
rect 9228 185 11300 194
rect 7276 151 7293 185
rect 7327 151 7465 185
rect 7499 151 7637 185
rect 7671 151 7809 185
rect 7843 151 7981 185
rect 8015 151 8153 185
rect 8187 151 8325 185
rect 8359 151 8497 185
rect 8531 151 8669 185
rect 8703 151 8841 185
rect 8875 151 9013 185
rect 9047 151 9176 185
rect 9228 151 9357 185
rect 9391 151 9529 185
rect 9563 151 9701 185
rect 9735 151 9873 185
rect 9907 151 10045 185
rect 10079 151 10217 185
rect 10251 151 10389 185
rect 10423 151 10561 185
rect 10595 151 10733 185
rect 10767 151 10905 185
rect 10939 151 11077 185
rect 11111 151 11249 185
rect 11283 151 11300 185
rect 7276 142 9176 151
rect 9228 142 11300 151
rect 7276 140 11300 142
<< via1 >>
rect 1264 4006 1316 4058
rect 2984 4006 3036 4058
rect 6854 4006 6906 4058
rect 9176 4006 9228 4058
rect 5478 3670 5530 3722
rect 6854 3670 6906 3722
rect 9176 3670 9228 3722
rect 1178 3629 1230 3638
rect 1178 3595 1187 3629
rect 1187 3595 1221 3629
rect 1221 3595 1230 3629
rect 1178 3586 1230 3595
rect 3070 3629 3122 3638
rect 3070 3595 3079 3629
rect 3079 3595 3113 3629
rect 3113 3595 3122 3629
rect 3070 3586 3122 3595
rect 6596 3586 6648 3638
rect 9262 3629 9314 3638
rect 9262 3595 9271 3629
rect 9271 3595 9305 3629
rect 9305 3595 9314 3629
rect 9262 3586 9314 3595
rect 4532 3250 4584 3302
rect 5478 3250 5530 3302
rect 1264 2914 1316 2966
rect 2984 2914 3036 2966
rect 4532 2914 4584 2966
rect 1264 2873 1316 2882
rect 1264 2839 1273 2873
rect 1273 2839 1307 2873
rect 1307 2839 1316 2873
rect 1264 2830 1316 2839
rect 2984 2873 3036 2882
rect 2984 2839 2993 2873
rect 2993 2839 3027 2873
rect 3027 2839 3036 2873
rect 2984 2830 3036 2839
rect 4274 2830 4326 2882
rect 5650 2830 5702 2882
rect 6854 2873 6906 2882
rect 6854 2839 6863 2873
rect 6863 2839 6897 2873
rect 6897 2839 6906 2873
rect 6854 2830 6906 2839
rect 9176 2873 9228 2882
rect 9176 2839 9185 2873
rect 9185 2839 9219 2873
rect 9219 2839 9228 2873
rect 9176 2830 9228 2839
rect 1092 2746 1144 2798
rect 2898 2746 2950 2798
rect 3156 2746 3208 2798
rect 9348 2746 9400 2798
rect 1092 2621 1144 2630
rect 1092 2587 1101 2621
rect 1101 2587 1135 2621
rect 1135 2587 1144 2621
rect 1092 2578 1144 2587
rect 3156 2621 3208 2630
rect 3156 2587 3165 2621
rect 3165 2587 3199 2621
rect 3199 2587 3208 2621
rect 3156 2578 3208 2587
rect 9348 2621 9400 2630
rect 9348 2587 9357 2621
rect 9357 2587 9391 2621
rect 9391 2587 9400 2621
rect 9348 2578 9400 2587
rect 1264 2494 1316 2546
rect 2984 2494 3036 2546
rect 5650 2494 5702 2546
rect 6854 2537 6906 2546
rect 6854 2503 6863 2537
rect 6863 2503 6897 2537
rect 6897 2503 6906 2537
rect 6854 2494 6906 2503
rect 9176 2494 9228 2546
rect 9348 2410 9400 2462
rect 4532 2158 4584 2210
rect 5478 2158 5530 2210
rect 4532 2117 4584 2126
rect 4532 2083 4541 2117
rect 4541 2083 4575 2117
rect 4575 2083 4584 2117
rect 4532 2074 4584 2083
rect 5478 2117 5530 2126
rect 5478 2083 5487 2117
rect 5487 2083 5521 2117
rect 5521 2083 5530 2117
rect 5478 2074 5530 2083
rect 4360 1990 4412 2042
rect 5564 2033 5616 2042
rect 5564 1999 5573 2033
rect 5573 1999 5607 2033
rect 5607 1999 5616 2033
rect 5564 1990 5616 1999
rect 4274 1906 4326 1958
rect 3070 1822 3122 1874
rect 4360 1865 4412 1874
rect 4360 1831 4369 1865
rect 4369 1831 4403 1865
rect 4403 1831 4412 1865
rect 4360 1822 4412 1831
rect 5564 1865 5616 1874
rect 5564 1831 5573 1865
rect 5573 1831 5607 1865
rect 5607 1831 5616 1865
rect 5564 1822 5616 1831
rect 1178 1738 1230 1790
rect 3070 1738 3122 1790
rect 4532 1738 4584 1790
rect 5478 1781 5530 1790
rect 5478 1747 5487 1781
rect 5487 1747 5521 1781
rect 5521 1747 5530 1781
rect 5478 1738 5530 1747
rect 6596 1738 6648 1790
rect 9262 1738 9314 1790
rect 1178 1486 1230 1538
rect 3156 1486 3208 1538
rect 1092 1445 1144 1454
rect 1092 1411 1101 1445
rect 1101 1411 1135 1445
rect 1135 1411 1144 1445
rect 1092 1402 1144 1411
rect 3156 1445 3208 1454
rect 3156 1411 3165 1445
rect 3165 1411 3199 1445
rect 3199 1411 3208 1445
rect 3156 1402 3208 1411
rect 9348 1445 9400 1454
rect 9348 1411 9357 1445
rect 9357 1411 9391 1445
rect 9391 1411 9400 1445
rect 9348 1402 9400 1411
rect 1264 1318 1316 1370
rect 2984 1318 3036 1370
rect 6854 1318 6906 1370
rect 9176 1318 9228 1370
rect 4274 982 4326 1034
rect 5650 982 5702 1034
rect 5478 898 5530 950
rect 6854 898 6906 950
rect 9176 898 9228 950
rect 2984 646 3036 698
rect 4532 646 4584 698
rect 5478 646 5530 698
rect 1178 562 1230 614
rect 3070 562 3122 614
rect 4532 605 4584 614
rect 4532 571 4541 605
rect 4541 571 4575 605
rect 4575 571 4584 605
rect 4532 562 4584 571
rect 5478 562 5530 614
rect 9262 562 9314 614
rect 1264 226 1316 278
rect 2984 226 3036 278
rect 1264 185 1316 194
rect 1264 151 1273 185
rect 1273 151 1307 185
rect 1307 151 1316 185
rect 1264 142 1316 151
rect 2984 185 3036 194
rect 2984 151 2993 185
rect 2993 151 3027 185
rect 3027 151 3036 185
rect 2984 142 3036 151
rect 9176 185 9228 194
rect 9176 151 9185 185
rect 9185 151 9219 185
rect 9219 151 9228 185
rect 9176 142 9228 151
<< metal2 >>
rect 1262 4058 1318 4064
rect 1262 4006 1264 4058
rect 1316 4006 1318 4058
rect 1176 3638 1232 3644
rect 1176 3586 1178 3638
rect 1230 3586 1232 3638
rect 1090 2798 1146 2804
rect 1090 2746 1092 2798
rect 1144 2746 1146 2798
rect 1090 2630 1146 2746
rect 1090 2578 1092 2630
rect 1144 2578 1146 2630
rect 1090 1454 1146 2578
rect 1090 1402 1092 1454
rect 1144 1402 1146 1454
rect 1090 1396 1146 1402
rect 1176 1790 1232 3586
rect 1262 2966 1318 4006
rect 1262 2914 1264 2966
rect 1316 2914 1318 2966
rect 1262 2882 1318 2914
rect 1262 2830 1264 2882
rect 1316 2830 1318 2882
rect 1262 2824 1318 2830
rect 2982 4058 3038 4064
rect 2982 4006 2984 4058
rect 3036 4006 3038 4058
rect 2982 2966 3038 4006
rect 6852 4058 6908 4064
rect 6852 4006 6854 4058
rect 6906 4006 6908 4058
rect 5476 3722 5532 3728
rect 5476 3670 5478 3722
rect 5530 3670 5532 3722
rect 2982 2914 2984 2966
rect 3036 2914 3038 2966
rect 2982 2882 3038 2914
rect 2982 2830 2984 2882
rect 3036 2830 3038 2882
rect 2982 2824 3038 2830
rect 3068 3638 3124 3644
rect 3068 3586 3070 3638
rect 3122 3586 3124 3638
rect 2896 2800 2952 2809
rect 2896 2735 2952 2744
rect 1176 1738 1178 1790
rect 1230 1738 1232 1790
rect 1176 1538 1232 1738
rect 1176 1486 1178 1538
rect 1230 1486 1232 1538
rect 1176 614 1232 1486
rect 1176 562 1178 614
rect 1230 562 1232 614
rect 1176 556 1232 562
rect 1262 2546 1318 2552
rect 1262 2494 1264 2546
rect 1316 2494 1318 2546
rect 1262 1370 1318 2494
rect 1262 1318 1264 1370
rect 1316 1318 1318 1370
rect 1262 278 1318 1318
rect 1262 226 1264 278
rect 1316 226 1318 278
rect 1262 194 1318 226
rect 1262 142 1264 194
rect 1316 142 1318 194
rect 1262 136 1318 142
rect 2982 2546 3038 2552
rect 2982 2494 2984 2546
rect 3036 2494 3038 2546
rect 2982 1370 3038 2494
rect 2982 1318 2984 1370
rect 3036 1318 3038 1370
rect 2982 698 3038 1318
rect 2982 646 2984 698
rect 3036 646 3038 698
rect 2982 278 3038 646
rect 3068 1874 3124 3586
rect 4530 3302 4586 3308
rect 4530 3250 4532 3302
rect 4584 3250 4586 3302
rect 4530 2966 4586 3250
rect 4530 2914 4532 2966
rect 4584 2914 4586 2966
rect 4272 2882 4328 2888
rect 4272 2830 4274 2882
rect 4326 2830 4328 2882
rect 3068 1822 3070 1874
rect 3122 1822 3124 1874
rect 3068 1790 3124 1822
rect 3068 1738 3070 1790
rect 3122 1738 3124 1790
rect 3068 614 3124 1738
rect 3154 2798 3210 2804
rect 3154 2746 3156 2798
rect 3208 2746 3210 2798
rect 3154 2630 3210 2746
rect 3154 2578 3156 2630
rect 3208 2578 3210 2630
rect 3154 1538 3210 2578
rect 3154 1486 3156 1538
rect 3208 1486 3210 1538
rect 3154 1454 3210 1486
rect 3154 1402 3156 1454
rect 3208 1402 3210 1454
rect 3154 1396 3210 1402
rect 4272 1958 4328 2830
rect 4530 2210 4586 2914
rect 4530 2158 4532 2210
rect 4584 2158 4586 2210
rect 4530 2126 4586 2158
rect 4530 2074 4532 2126
rect 4584 2074 4586 2126
rect 4530 2068 4586 2074
rect 5476 3302 5532 3670
rect 6852 3722 6908 4006
rect 6852 3670 6854 3722
rect 6906 3670 6908 3722
rect 5476 3250 5478 3302
rect 5530 3250 5532 3302
rect 5476 2210 5532 3250
rect 6594 3638 6650 3644
rect 6594 3586 6596 3638
rect 6648 3586 6650 3638
rect 5476 2158 5478 2210
rect 5530 2158 5532 2210
rect 5476 2126 5532 2158
rect 5476 2074 5478 2126
rect 5530 2074 5532 2126
rect 5476 2068 5532 2074
rect 5648 2882 5704 2888
rect 5648 2830 5650 2882
rect 5702 2830 5704 2882
rect 5648 2546 5704 2830
rect 5648 2494 5650 2546
rect 5702 2494 5704 2546
rect 4272 1906 4274 1958
rect 4326 1906 4328 1958
rect 4272 1034 4328 1906
rect 4358 2042 4414 2048
rect 4358 1990 4360 2042
rect 4412 1990 4414 2042
rect 4358 1874 4414 1990
rect 4358 1822 4360 1874
rect 4412 1822 4414 1874
rect 4358 1816 4414 1822
rect 5562 2042 5618 2048
rect 5562 1990 5564 2042
rect 5616 1990 5618 2042
rect 5562 1874 5618 1990
rect 5562 1822 5564 1874
rect 5616 1822 5618 1874
rect 5562 1816 5618 1822
rect 4272 982 4274 1034
rect 4326 982 4328 1034
rect 4272 976 4328 982
rect 4530 1790 4586 1796
rect 4530 1738 4532 1790
rect 4584 1738 4586 1790
rect 3068 562 3070 614
rect 3122 562 3124 614
rect 3068 556 3124 562
rect 4530 698 4586 1738
rect 4530 646 4532 698
rect 4584 646 4586 698
rect 4530 614 4586 646
rect 4530 562 4532 614
rect 4584 562 4586 614
rect 4530 556 4586 562
rect 5476 1790 5532 1796
rect 5476 1738 5478 1790
rect 5530 1738 5532 1790
rect 5476 950 5532 1738
rect 5648 1034 5704 2494
rect 6594 1790 6650 3586
rect 6852 2882 6908 3670
rect 6852 2830 6854 2882
rect 6906 2830 6908 2882
rect 6852 2824 6908 2830
rect 9174 4058 9230 4064
rect 9174 4006 9176 4058
rect 9228 4006 9230 4058
rect 9174 3722 9230 4006
rect 9174 3670 9176 3722
rect 9228 3670 9230 3722
rect 9174 2882 9230 3670
rect 9174 2830 9176 2882
rect 9228 2830 9230 2882
rect 9174 2824 9230 2830
rect 9260 3638 9316 3644
rect 9260 3586 9262 3638
rect 9314 3586 9316 3638
rect 9260 2800 9316 3586
rect 6594 1738 6596 1790
rect 6648 1738 6650 1790
rect 6594 1732 6650 1738
rect 6852 2546 6908 2552
rect 6852 2494 6854 2546
rect 6906 2494 6908 2546
rect 5648 982 5650 1034
rect 5702 982 5704 1034
rect 5648 976 5704 982
rect 6852 1370 6908 2494
rect 6852 1318 6854 1370
rect 6906 1318 6908 1370
rect 5476 898 5478 950
rect 5530 898 5532 950
rect 5476 698 5532 898
rect 6852 950 6908 1318
rect 6852 898 6854 950
rect 6906 898 6908 950
rect 6852 892 6908 898
rect 9174 2546 9230 2552
rect 9174 2494 9176 2546
rect 9228 2494 9230 2546
rect 9174 1370 9230 2494
rect 9174 1318 9176 1370
rect 9228 1318 9230 1370
rect 9174 950 9230 1318
rect 9174 898 9176 950
rect 9228 898 9230 950
rect 5476 646 5478 698
rect 5530 646 5532 698
rect 5476 614 5532 646
rect 5476 562 5478 614
rect 5530 562 5532 614
rect 5476 556 5532 562
rect 2982 226 2984 278
rect 3036 226 3038 278
rect 2982 194 3038 226
rect 2982 142 2984 194
rect 3036 142 3038 194
rect 2982 136 3038 142
rect 9174 194 9230 898
rect 9260 1790 9316 2744
rect 9260 1738 9262 1790
rect 9314 1738 9316 1790
rect 9260 614 9316 1738
rect 9346 2798 9402 2804
rect 9346 2746 9348 2798
rect 9400 2746 9402 2798
rect 9346 2630 9402 2746
rect 9346 2578 9348 2630
rect 9400 2578 9402 2630
rect 9346 2462 9402 2578
rect 9346 2410 9348 2462
rect 9400 2410 9402 2462
rect 9346 1454 9402 2410
rect 9346 1402 9348 1454
rect 9400 1402 9402 1454
rect 9346 1396 9402 1402
rect 9260 562 9262 614
rect 9314 562 9316 614
rect 9260 556 9316 562
rect 9174 142 9176 194
rect 9228 142 9230 194
rect 9174 136 9230 142
<< via2 >>
rect 2896 2798 2952 2800
rect 2896 2746 2898 2798
rect 2898 2746 2950 2798
rect 2950 2746 2952 2798
rect 2896 2744 2952 2746
rect 9260 2744 9316 2800
<< metal3 >>
rect 2891 2800 9321 2852
rect 2891 2744 2896 2800
rect 2952 2744 9260 2800
rect 9316 2744 9321 2800
rect 2891 2692 9321 2744
<< labels >>
flabel locali 7285 2210 7335 2587 0 FreeSans 1600 0 0 0 clkout
port 0 nsew
flabel poly 6220 1092 6250 1302 0 FreeSans 1600 0 0 0 clk1
port 1 nsew
flabel pwell 6751 3894 6837 4170 0 FreeSans 1600 0 0 0 gnd
port 2 nsew
flabel nwell 6536 1176 11524 2688 0 FreeSans 1600 0 0 0 vdd
port 4 nsew
<< end >>
