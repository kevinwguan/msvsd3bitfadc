MACRO INV_80711309
  ORIGIN 0 0 ;
  FOREIGN INV_80711309 0 0 ;
  SIZE 22.36 BY 21 ;
  PIN ZN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 11.47 7.82 11.75 14.02 ;
      LAYER M2 ;
        RECT 11.01 7 12.21 7.28 ;
      LAYER M3 ;
        RECT 11.47 7.14 11.75 7.98 ;
      LAYER M2 ;
        RECT 11.45 7 11.77 7.28 ;
    END
  END ZN
  PIN I
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 11.04 12.02 11.32 18.22 ;
      LAYER M2 ;
        RECT 11.01 2.8 12.21 3.08 ;
      LAYER M3 ;
        RECT 11.04 2.94 11.32 12.18 ;
      LAYER M2 ;
        RECT 11.02 2.8 11.34 3.08 ;
    END
  END I
  PIN SN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 10.61 0.68 10.89 6.88 ;
    END
  END SN
  PIN SP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 10.61 8.24 10.89 20.32 ;
    END
  END SP
  OBS 
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 11.055 2.435 11.305 3.445 ;
  LAYER M1 ;
        RECT 11.055 0.335 11.305 1.345 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M2 ;
        RECT 10.58 6.58 11.78 6.86 ;
  LAYER M2 ;
        RECT 10.58 0.7 11.78 0.98 ;
  LAYER M2 ;
        RECT 11.01 7 12.21 7.28 ;
  LAYER M2 ;
        RECT 11.01 2.8 12.21 3.08 ;
  LAYER M3 ;
        RECT 10.61 0.68 10.89 6.88 ;
  LAYER M1 ;
        RECT 20.945 7.895 21.195 11.425 ;
  LAYER M1 ;
        RECT 20.945 11.675 21.195 12.685 ;
  LAYER M1 ;
        RECT 20.945 13.775 21.195 17.305 ;
  LAYER M1 ;
        RECT 20.945 17.555 21.195 18.565 ;
  LAYER M1 ;
        RECT 20.945 19.655 21.195 20.665 ;
  LAYER M1 ;
        RECT 21.375 7.895 21.625 11.425 ;
  LAYER M1 ;
        RECT 21.375 13.775 21.625 17.305 ;
  LAYER M1 ;
        RECT 20.515 7.895 20.765 11.425 ;
  LAYER M1 ;
        RECT 20.515 13.775 20.765 17.305 ;
  LAYER M1 ;
        RECT 20.085 7.895 20.335 11.425 ;
  LAYER M1 ;
        RECT 20.085 11.675 20.335 12.685 ;
  LAYER M1 ;
        RECT 20.085 13.775 20.335 17.305 ;
  LAYER M1 ;
        RECT 20.085 17.555 20.335 18.565 ;
  LAYER M1 ;
        RECT 20.085 19.655 20.335 20.665 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M1 ;
        RECT 19.655 13.775 19.905 17.305 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 11.425 ;
  LAYER M1 ;
        RECT 19.225 11.675 19.475 12.685 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 17.305 ;
  LAYER M1 ;
        RECT 19.225 17.555 19.475 18.565 ;
  LAYER M1 ;
        RECT 19.225 19.655 19.475 20.665 ;
  LAYER M1 ;
        RECT 18.795 7.895 19.045 11.425 ;
  LAYER M1 ;
        RECT 18.795 13.775 19.045 17.305 ;
  LAYER M1 ;
        RECT 18.365 7.895 18.615 11.425 ;
  LAYER M1 ;
        RECT 18.365 11.675 18.615 12.685 ;
  LAYER M1 ;
        RECT 18.365 13.775 18.615 17.305 ;
  LAYER M1 ;
        RECT 18.365 17.555 18.615 18.565 ;
  LAYER M1 ;
        RECT 18.365 19.655 18.615 20.665 ;
  LAYER M1 ;
        RECT 17.935 7.895 18.185 11.425 ;
  LAYER M1 ;
        RECT 17.935 13.775 18.185 17.305 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 11.425 ;
  LAYER M1 ;
        RECT 17.505 11.675 17.755 12.685 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 17.305 ;
  LAYER M1 ;
        RECT 17.505 17.555 17.755 18.565 ;
  LAYER M1 ;
        RECT 17.505 19.655 17.755 20.665 ;
  LAYER M1 ;
        RECT 17.075 7.895 17.325 11.425 ;
  LAYER M1 ;
        RECT 17.075 13.775 17.325 17.305 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 11.425 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 12.685 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 17.305 ;
  LAYER M1 ;
        RECT 16.645 17.555 16.895 18.565 ;
  LAYER M1 ;
        RECT 16.645 19.655 16.895 20.665 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M1 ;
        RECT 16.215 13.775 16.465 17.305 ;
  LAYER M1 ;
        RECT 15.785 7.895 16.035 11.425 ;
  LAYER M1 ;
        RECT 15.785 11.675 16.035 12.685 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 17.305 ;
  LAYER M1 ;
        RECT 15.785 17.555 16.035 18.565 ;
  LAYER M1 ;
        RECT 15.785 19.655 16.035 20.665 ;
  LAYER M1 ;
        RECT 15.355 7.895 15.605 11.425 ;
  LAYER M1 ;
        RECT 15.355 13.775 15.605 17.305 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 11.425 ;
  LAYER M1 ;
        RECT 14.925 11.675 15.175 12.685 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 17.305 ;
  LAYER M1 ;
        RECT 14.925 17.555 15.175 18.565 ;
  LAYER M1 ;
        RECT 14.925 19.655 15.175 20.665 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 14.495 13.775 14.745 17.305 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 17.305 ;
  LAYER M1 ;
        RECT 14.065 17.555 14.315 18.565 ;
  LAYER M1 ;
        RECT 14.065 19.655 14.315 20.665 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 13.635 13.775 13.885 17.305 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 11.425 ;
  LAYER M1 ;
        RECT 13.205 11.675 13.455 12.685 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 17.305 ;
  LAYER M1 ;
        RECT 13.205 17.555 13.455 18.565 ;
  LAYER M1 ;
        RECT 13.205 19.655 13.455 20.665 ;
  LAYER M1 ;
        RECT 12.775 7.895 13.025 11.425 ;
  LAYER M1 ;
        RECT 12.775 13.775 13.025 17.305 ;
  LAYER M1 ;
        RECT 12.345 7.895 12.595 11.425 ;
  LAYER M1 ;
        RECT 12.345 11.675 12.595 12.685 ;
  LAYER M1 ;
        RECT 12.345 13.775 12.595 17.305 ;
  LAYER M1 ;
        RECT 12.345 17.555 12.595 18.565 ;
  LAYER M1 ;
        RECT 12.345 19.655 12.595 20.665 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M1 ;
        RECT 11.915 13.775 12.165 17.305 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 17.305 ;
  LAYER M1 ;
        RECT 11.485 17.555 11.735 18.565 ;
  LAYER M1 ;
        RECT 11.485 19.655 11.735 20.665 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M1 ;
        RECT 11.055 13.775 11.305 17.305 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 11.425 ;
  LAYER M1 ;
        RECT 10.625 11.675 10.875 12.685 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 17.305 ;
  LAYER M1 ;
        RECT 10.625 17.555 10.875 18.565 ;
  LAYER M1 ;
        RECT 10.625 19.655 10.875 20.665 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 10.195 13.775 10.445 17.305 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 17.305 ;
  LAYER M1 ;
        RECT 9.765 17.555 10.015 18.565 ;
  LAYER M1 ;
        RECT 9.765 19.655 10.015 20.665 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 9.335 13.775 9.585 17.305 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 17.305 ;
  LAYER M1 ;
        RECT 8.905 17.555 9.155 18.565 ;
  LAYER M1 ;
        RECT 8.905 19.655 9.155 20.665 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 8.475 13.775 8.725 17.305 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 17.305 ;
  LAYER M1 ;
        RECT 8.045 17.555 8.295 18.565 ;
  LAYER M1 ;
        RECT 8.045 19.655 8.295 20.665 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M1 ;
        RECT 7.615 13.775 7.865 17.305 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 11.425 ;
  LAYER M1 ;
        RECT 7.185 11.675 7.435 12.685 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 17.305 ;
  LAYER M1 ;
        RECT 7.185 17.555 7.435 18.565 ;
  LAYER M1 ;
        RECT 7.185 19.655 7.435 20.665 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 6.755 13.775 7.005 17.305 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 17.305 ;
  LAYER M1 ;
        RECT 6.325 17.555 6.575 18.565 ;
  LAYER M1 ;
        RECT 6.325 19.655 6.575 20.665 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M1 ;
        RECT 5.895 13.775 6.145 17.305 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 11.425 ;
  LAYER M1 ;
        RECT 5.465 11.675 5.715 12.685 ;
  LAYER M1 ;
        RECT 5.465 13.775 5.715 17.305 ;
  LAYER M1 ;
        RECT 5.465 17.555 5.715 18.565 ;
  LAYER M1 ;
        RECT 5.465 19.655 5.715 20.665 ;
  LAYER M1 ;
        RECT 5.035 7.895 5.285 11.425 ;
  LAYER M1 ;
        RECT 5.035 13.775 5.285 17.305 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 11.425 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 12.685 ;
  LAYER M1 ;
        RECT 4.605 13.775 4.855 17.305 ;
  LAYER M1 ;
        RECT 4.605 17.555 4.855 18.565 ;
  LAYER M1 ;
        RECT 4.605 19.655 4.855 20.665 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 4.175 13.775 4.425 17.305 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 17.305 ;
  LAYER M1 ;
        RECT 3.745 17.555 3.995 18.565 ;
  LAYER M1 ;
        RECT 3.745 19.655 3.995 20.665 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 3.315 13.775 3.565 17.305 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 11.425 ;
  LAYER M1 ;
        RECT 2.885 11.675 3.135 12.685 ;
  LAYER M1 ;
        RECT 2.885 13.775 3.135 17.305 ;
  LAYER M1 ;
        RECT 2.885 17.555 3.135 18.565 ;
  LAYER M1 ;
        RECT 2.885 19.655 3.135 20.665 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 2.455 13.775 2.705 17.305 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 17.305 ;
  LAYER M1 ;
        RECT 2.025 17.555 2.275 18.565 ;
  LAYER M1 ;
        RECT 2.025 19.655 2.275 20.665 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 1.595 13.775 1.845 17.305 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 17.305 ;
  LAYER M1 ;
        RECT 1.165 17.555 1.415 18.565 ;
  LAYER M1 ;
        RECT 1.165 19.655 1.415 20.665 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 0.735 13.775 0.985 17.305 ;
  LAYER M2 ;
        RECT 1.12 7.84 21.24 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 21.24 12.32 ;
  LAYER M2 ;
        RECT 0.69 8.26 21.67 8.54 ;
  LAYER M2 ;
        RECT 1.12 13.72 21.24 14 ;
  LAYER M2 ;
        RECT 1.12 17.92 21.24 18.2 ;
  LAYER M2 ;
        RECT 0.69 14.14 21.67 14.42 ;
  LAYER M2 ;
        RECT 1.12 20.02 21.24 20.3 ;
  LAYER M3 ;
        RECT 11.47 7.82 11.75 14.02 ;
  LAYER M3 ;
        RECT 11.04 12.02 11.32 18.22 ;
  LAYER M3 ;
        RECT 10.61 8.24 10.89 20.32 ;
  END 
END INV_80711309
